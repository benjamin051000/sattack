//# 35 inputs
//# 49 outputs
//# 179 D-type flipflops
//# 1775 inverters
//# 1004 gates (0 ANDs + 0 NANDs + 239 ORs + 765 NORs)

module dff (CK,Q,D);
input CK,D;
output Q;

  always @(posedge CK)
    Q <= D;

endmodule

module s5378(GND,VDD,CK,n3065gat,n3066gat,n3067gat,n3068gat,n3069gat,n3070gat,
n3071gat,
n3072gat,n3073gat,n3074gat,n3075gat,n3076gat,n3077gat,n3078gat,n3079gat,
n3080gat,n3081gat,n3082gat,n3083gat,n3084gat,n3085gat,n3086gat,n3087gat,
n3088gat,n3089gat,n3090gat,n3091gat,n3092gat,n3093gat,n3094gat,n3095gat,
n3097gat,n3098gat,n3099gat,n3100gat,n3104gat,n3105gat,n3106gat,n3107gat,
n3108gat,n3109gat,n3110gat,n3111gat,n3112gat,n3113gat,n3114gat,n3115gat,
n3116gat,n3117gat,n3118gat,n3119gat,n3120gat,n3121gat,n3122gat,n3123gat,
n3124gat,n3125gat,n3126gat,n3127gat,n3128gat,n3129gat,n3130gat,n3131gat,
n3132gat,n3133gat,n3134gat,n3135gat,n3136gat,n3137gat,n3138gat,n3139gat,
n3140gat,n3141gat,n3142gat,n3143gat,n3144gat,n3145gat,n3146gat,n3147gat,
n3148gat,n3149gat,n3150gat,n3151gat,n3152gat);
input GND,VDD,CK,n3065gat,n3066gat,n3067gat,n3068gat,n3069gat,n3070gat,
n3071gat,n3072gat,
n3073gat,n3074gat,n3075gat,n3076gat,n3077gat,n3078gat,n3079gat,n3080gat,
n3081gat,n3082gat,n3083gat,n3084gat,n3085gat,n3086gat,n3087gat,n3088gat,
n3089gat,n3090gat,n3091gat,n3092gat,n3093gat,n3094gat,n3095gat,n3097gat,
n3098gat,n3099gat,n3100gat;
output n3104gat,n3105gat,n3106gat,n3107gat,n3108gat,n3109gat,n3110gat,n3111gat,
n3112gat,n3113gat,n3114gat,n3115gat,n3116gat,n3117gat,n3118gat,n3119gat,
n3120gat,n3121gat,n3122gat,n3123gat,n3124gat,n3125gat,n3126gat,n3127gat,
n3128gat,n3129gat,n3130gat,n3131gat,n3132gat,n3133gat,n3134gat,n3135gat,
n3136gat,n3137gat,n3138gat,n3139gat,n3140gat,n3141gat,n3142gat,n3143gat,
n3144gat,n3145gat,n3146gat,n3147gat,n3148gat,n3149gat,n3150gat,n3151gat,
n3152gat;

wire n673gat,n2897gat,n398gat,n2782gat,n402gat,n2790gat,n919gat,n2670gat,
  n846gat,n2793gat,n394gat,n703gat,n722gat,n726gat,n2510gat,n748gat,n271gat,
  n2732gat,n160gat,n2776gat,n337gat,n2735gat,n842gat,n2673gat,n341gat,
  n2779gat,n2522gat,n43gat,n2472gat,n1620gat,n2319gat,n2470gat,n1821gat,
  n1827gat,n1825gat,n2029gat,n1816gat,n1829gat,n2027gat,n283gat,n165gat,
  n279gat,n1026gat,n275gat,n2476gat,n55gat,n1068gat,n2914gat,n957gat,
  n2928gat,n861gat,n2927gat,n1294gat,n2896gat,n1241gat,n2922gat,n1298gat,
  n865gat,n2894gat,n1080gat,n2921gat,n1148gat,n2895gat,n2468gat,n933gat,
  n618gat,n491gat,n622gat,n626gat,n834gat,n3064gat,n707gat,n3055gat,n838gat,
  n3063gat,n830gat,n3062gat,n614gat,n3056gat,n2526gat,n504gat,n680gat,
  n2913gat,n816gat,n2920gat,n580gat,n2905gat,n824gat,n3057gat,n820gat,
  n3059gat,n883gat,n3058gat,n584gat,n2898gat,n684gat,n3060gat,n699gat,
  n3061gat,n2464gat,n567gat,n2399gat,n3048gat,n2343gat,n3049gat,n2203gat,
  n3051gat,n2562gat,n3047gat,n2207gat,n3050gat,n2626gat,n3040gat,n2490gat,
  n3044gat,n2622gat,n3042gat,n2630gat,n3037gat,n2543gat,n3041gat,n2102gat,
  n1606gat,n1880gat,n3052gat,n1763gat,n1610gat,n2155gat,n1858gat,n1035gat,
  n2918gat,n1121gat,n2952gat,n1072gat,n2919gat,n1282gat,n2910gat,n1226gat,
  n2907gat,n931gat,n2911gat,n1135gat,n2912gat,n1045gat,n2909gat,n1197gat,
  n2908gat,n2518gat,n2971gat,n667gat,n2904gat,n659gat,n2891gat,n553gat,
  n2903gat,n777gat,n2915gat,n561gat,n2901gat,n366gat,n2890gat,n322gat,
  n2888gat,n318gat,n2887gat,n314gat,n2886gat,n2599gat,n3010gat,n2588gat,
  n3016gat,n2640gat,n3054gat,n2658gat,n2579gat,n2495gat,n3036gat,n2390gat,
  n3034gat,n2270gat,n3031gat,n2339gat,n3035gat,n2502gat,n2646gat,n2634gat,
  n3053gat,n2506gat,n2613gat,n1834gat,n1625gat,n1767gat,n1626gat,n2084gat,
  n1603gat,n2143gat,n2541gat,n2061gat,n2557gat,n2139gat,n2487gat,n1899gat,
  n2532gat,n1850gat,n2628gat,n2403gat,n2397gat,n2394gat,n2341gat,n2440gat,
  n2560gat,n2407gat,n2205gat,n2347gat,n2201gat,n1389gat,n1793gat,n2021gat,
  n1781gat,n1394gat,n1516gat,n1496gat,n1392gat,n2091gat,n1685gat,n1332gat,
  n1565gat,n1740gat,n1330gat,n2179gat,n1945gat,n2190gat,n2268gat,n2135gat,
  n2337gat,n2262gat,n2388gat,n2182gat,n1836gat,n1433gat,n2983gat,n1316gat,
  n1431gat,n1363gat,n1314gat,n1312gat,n1361gat,n1775gat,n1696gat,n1871gat,
  n2009gat,n2592gat,n1773gat,n1508gat,n1636gat,n1678gat,n1712gat,n2309gat,
  n3000gat,n2450gat,n2307gat,n2446gat,n2661gat,n2095gat,n827gat,n2176gat,
  n2093gat,n2169gat,n2174gat,n2454gat,n2163gat,n2040gat,n1777gat,n2044gat,
  n2015gat,n2037gat,n2042gat,n2025gat,n2017gat,n2099gat,n2023gat,n2266gat,
  n2493gat,n2033gat,n2035gat,n2110gat,n2031gat,n2125gat,n2108gat,n2121gat,
  n2123gat,n2117gat,n2119gat,n1975gat,n2632gat,n2644gat,n2638gat,n156gat,
  n612gat,n152gat,n705gat,n331gat,n822gat,n388gat,n881gat,n463gat,n818gat,
  n327gat,n682gat,n384gat,n697gat,n256gat,n836gat,n470gat,n828gat,n148gat,
  n832gat,n2458gat,n2590gat,n2514gat,n2456gat,n1771gat,n1613gat,n1336gat,
  n1391gat,n1748gat,n1927gat,n1675gat,n1713gat,n1807gat,n1717gat,n1340gat,
  n1567gat,n1456gat,n1564gat,n1525gat,n1632gat,n1462gat,n1915gat,n1596gat,
  n1800gat,n1588gat,n1593gat,II1,n2717gat,n2715gat,II5,n2725gat,n2723gat,
  n296gat,n421gat,II11,n2768gat,II14,n2767gat,n373gat,II18,n2671gat,n2669gat,
  II23,n2845gat,n2844gat,II27,n2668gat,II30,n2667gat,n856gat,II44,n672gat,
  II47,n2783gat,II50,n396gat,II62,n2791gat,II65,II76,n401gat,n1645gat,
  n1499gat,II81,II92,n918gat,n1553gat,n1616gat,II97,n2794gat,II100,II111,
  n845gat,n1559gat,n1614gat,n1643gat,n1641gat,n1651gat,n1642gat,n1562gat,
  n1556gat,n1560gat,n1557gat,n1640gat,n1639gat,n1566gat,n1605gat,n1554gat,
  n1555gat,n1722gat,n1558gat,n392gat,II149,n702gat,n1319gat,n1256gat,n720gat,
  II171,n725gat,n1447gat,n1117gat,n1627gat,n1618gat,II178,n721gat,n1380gat,
  n1114gat,n1628gat,n1621gat,n701gat,n1446gat,n1318gat,n1705gat,n1619gat,
  n1706gat,n1622gat,II192,n2856gat,n2854gat,II196,n1218gat,II199,n2861gat,
  n2859gat,II203,n1219gat,II206,n2864gat,n2862gat,II210,n1220gat,II214,
  n2860gat,II217,n1221gat,II220,n2863gat,II223,n1222gat,II227,n2855gat,II230,
  n1223gat,n640gat,n1213gat,II237,n753gat,II240,n2716gat,II243,n2869gat,
  n2867gat,II248,n2868gat,II253,n2906gat,n754gat,II256,n2724gat,II259,
  n2728gat,n2726gat,II264,n2727gat,n422gat,n2889gat,II270,n755gat,n747gat,
  II275,n756gat,II278,n757gat,II282,n758gat,n2508gat,II297,n2733gat,II300,
  II311,n270gat,II314,n263gat,II317,n2777gat,II320,II331,n159gat,II334,
  n264gat,II337,n2736gat,II340,II351,n336gat,II354,n265gat,n158gat,II359,
  n266gat,n335gat,II363,n267gat,n269gat,II368,n268gat,n41gat,n258gat,II375,
  n48gat,II378,n1018gat,II381,n2674gat,II384,II395,n841gat,II398,n1019gat,
  II401,n1020gat,n840gat,II406,n1021gat,II409,n1022gat,n724gat,II414,
  n1023gat,II420,n1013gat,n49gat,II423,n2780gat,II426,II437,n340gat,II440,
  n480gat,II443,n481gat,II446,n393gat,II449,n482gat,II453,n483gat,II456,
  n484gat,n339gat,II461,n485gat,n42gat,n475gat,II468,n50gat,n162gat,II473,
  n51gat,II476,n52gat,II480,n53gat,n2520gat,n1448gat,n1376gat,n1701gat,
  n1617gat,n1379gat,n1377gat,n1615gat,n1624gat,n1500gat,n1113gat,n1503gat,
  n1501gat,n1779gat,n1623gat,II509,n2730gat,II512,n2729gat,n2317gat,n1819gat,
  n1823gat,n1817gat,II572,n1828gat,II576,n2851gat,II579,n2850gat,II583,
  n2786gat,n2785gat,n92gat,n637gat,n529gat,n293gat,n361gat,II591,n2722gat,
  II594,n2721gat,n297gat,II606,n282gat,II609,n172gat,II620,n164gat,II623,
  n173gat,II634,n278gat,II637,n174gat,n163gat,II642,n175gat,n277gat,II646,
  n176gat,n281gat,II651,n177gat,n54gat,n167gat,II658,n60gat,II661,n911gat,
  II672,n1025gat,II675,n912gat,II678,n913gat,n1024gat,II683,n914gat,n917gat,
  II687,n915gat,n844gat,II692,n916gat,II698,n906gat,n61gat,II709,n274gat,
  II712,n348gat,II715,n349gat,II718,n397gat,II721,n350gat,n400gat,II726,
  n351gat,II729,n352gat,n273gat,II734,n353gat,n178gat,n343gat,II741,n62gat,
  n66gat,II746,n63gat,II749,n64gat,II753,n65gat,n2474gat,II768,n2832gat,
  II771,n2831gat,n2731gat,II776,n2719gat,n2718gat,II790,n1067gat,II793,
  n949gat,II796,n2839gat,n2838gat,n2775gat,II812,n956gat,II815,n950gat,II818,
  n2712gat,n2711gat,n2734gat,II834,n860gat,II837,n951gat,n955gat,II842,
  n952gat,n859gat,II846,n953gat,n1066gat,II851,n954gat,n857gat,n944gat,II858,
  n938gat,n2792gat,II863,n2847gat,n2846gat,II877,n1293gat,II880,n1233gat,
  n2672gat,II885,n2853gat,n2852gat,II899,n1240gat,II902,n1234gat,II913,
  n1297gat,II916,n1235gat,n1239gat,II921,n1236gat,n1296gat,II925,n1237gat,
  n1292gat,II930,n1238gat,II936,n1228gat,n939gat,n2778gat,II941,n2837gat,
  n2836gat,II955,n864gat,II958,n1055gat,n2789gat,II963,n2841gat,n2840gat,
  II977,n1079gat,II980,n1056gat,n2781gat,II985,n2843gat,n2842gat,II999,
  n1147gat,II1002,n1057gat,n1078gat,II1007,n1058gat,n1146gat,II1011,n1059gat,
  n863gat,II1016,n1060gat,n928gat,n1050gat,II1023,n940gat,n858gat,II1028,
  n941gat,II1031,n942gat,II1035,n943gat,n2466gat,n2720gat,n740gat,n2784gat,
  n743gat,n746gat,n294gat,n360gat,n374gat,n616gat,II1067,n501gat,n489gat,
  II1079,n502gat,II1082,n617gat,II1085,n499gat,II1088,n490gat,II1091,n500gat,
  n620gat,II1103,n738gat,n624gat,II1115,n737gat,II1118,n621gat,II1121,
  n733gat,II1124,n625gat,II1127,n735gat,II1138,n833gat,II1141,n714gat,II1152,
  n706gat,II1155,n715gat,II1166,n837gat,II1169,n716gat,II1174,n717gat,II1178,
  n718gat,II1183,n719gat,n515gat,n709gat,II1190,n509gat,II1201,n829gat,
  II1204,n734gat,II1209,n736gat,II1216,n728gat,n510gat,II1227,n613gat,II1230,
  n498gat,II1236,n503gat,n404gat,n493gat,II1243,n511gat,n405gat,II1248,
  n512gat,II1251,n513gat,II1255,n514gat,n2524gat,n17gat,n564gat,n79gat,
  n86gat,n219gat,n78gat,n563gat,II1278,n289gat,n179gat,n287gat,n188gat,
  n288gat,n72gat,n181gat,n111gat,n182gat,II1302,n679gat,II1305,n808gat,
  II1319,n815gat,II1322,n809gat,II1336,n579gat,II1339,n810gat,n814gat,II1344,
  n811gat,n578gat,II1348,n812gat,n678gat,II1353,n813gat,n677gat,n803gat,
  II1360,n572gat,II1371,n823gat,II1374,n591gat,II1385,n819gat,II1388,n592gat,
  II1399,n882gat,II1402,n593gat,II1407,n594gat,II1411,n595gat,II1416,n596gat,
  II1422,n586gat,n573gat,II1436,n583gat,II1439,n691gat,II1450,n683gat,II1453,
  n692gat,II1464,n698gat,II1467,n693gat,II1472,n694gat,II1476,n695gat,
  n582gat,II1481,n696gat,n456gat,n686gat,II1488,n574gat,n565gat,II1493,
  n575gat,II1496,n576gat,II1500,n577gat,n2462gat,n2665gat,II1516,n2596gat,
  n189gat,n286gat,n194gat,n187gat,n21gat,n15gat,II1538,n2398gat,n2353gat,
  II1550,n2342gat,n2284gat,n2354gat,n2356gat,n2214gat,n2286gat,II1585,
  n2624gat,II1606,n2489gat,II1617,n2621gat,n2533gat,n2534gat,II1630,n2629gat,
  n2486gat,n2429gat,n2432gat,n2430gat,II1655,n2101gat,n1693gat,II1667,
  n1879gat,n1698gat,n1934gat,n1543gat,II1683,n1762gat,n1673gat,n2989gat,
  II1698,n2154gat,n2488gat,II1703,n2625gat,n2530gat,n2531gat,II1708,n2542gat,
  n2482gat,n2426gat,n2480gat,n2153gat,n2355gat,II1719,n2561gat,n2443gat,
  n2289gat,II1724,n2148gat,II1734,n855gat,n759gat,II1749,n1034gat,II1752,
  n1189gat,n1075gat,II1766,n1120gat,II1769,n1190gat,n760gat,II1783,n1071gat,
  II1786,n1191gat,n1119gat,II1791,n1192gat,n1070gat,II1795,n1193gat,n1033gat,
  II1800,n1194gat,n1183gat,n1184gat,II1807,n1274gat,n644gat,n1280gat,n641gat,
  II1833,n1225gat,II1837,n1281gat,n1224gat,II1843,n2970gat,n1275gat,n761gat,
  II1857,n930gat,II1860,n1206gat,n762gat,II1874,n1134gat,II1877,n1207gat,
  n643gat,II1891,n1044gat,II1894,n1208gat,n1133gat,II1899,n1209gat,n1043gat,
  II1903,n1210gat,n929gat,II1908,n1211gat,n1268gat,n1201gat,II1915,n1276gat,
  n1329gat,II1920,n1277gat,II1923,n1278gat,II1927,n1279gat,n1284gat,n1269gat,
  n642gat,n1195gat,II1947,n1196gat,n2516gat,II1961,n3017gat,n851gat,n853gat,
  n1725gat,n664gat,n852gat,n854gat,II1981,n666gat,n368gat,II1996,n658gat,
  II1999,n784gat,n662gat,II2014,n552gat,II2017,n785gat,n661gat,II2032,
  n776gat,II2035,n786gat,n551gat,II2040,n787gat,n775gat,II2044,n788gat,
  n657gat,II2049,n789gat,n35gat,n779gat,II2056,n125gat,n558gat,n559gat,
  n371gat,II2084,n365gat,II2088,n560gat,n364gat,II2094,n2876gat,n126gat,
  n663gat,II2109,n321gat,II2112,n226gat,n370gat,II2127,n317gat,II2130,
  n227gat,n369gat,II2145,n313gat,II2148,n228gat,n316gat,II2153,n229gat,
  n312gat,II2157,n230gat,n320gat,II2162,n231gat,n34gat,n221gat,II2169,
  n127gat,n133gat,II2174,n128gat,II2177,n129gat,II2181,n130gat,n665gat,
  n1601gat,n120gat,n2597gat,n2595gat,n2594gat,n2586gat,II2213,n2573gat,
  II2225,n2574gat,II2228,n2575gat,II2232,n2639gat,II2235,n2576gat,II2238,
  n2577gat,II2242,n2578gat,II2248,n2568gat,n2582gat,II2251,n2206gat,II2254,
  n2414gat,II2257,n2415gat,II2260,n2202gat,II2263,n2416gat,II2268,n2417gat,
  II2271,n2418gat,II2275,n2419gat,II2281,n2409gat,n2585gat,n2656gat,II2316,
  n2389gat,II2319,n2494gat,II2324,n3014gat,n2649gat,II2344,n2338gat,II2349,
  n2269gat,II2354,n2880gat,n2652gat,n2500gat,n2620gat,n2612gat,II2372,
  n2606gat,II2376,n2607gat,n2540gat,II2380,n2608gat,n2536gat,II2385,n2609gat,
  II2389,n2610gat,II2394,n2611gat,II2400,n2601gat,n2616gat,II2403,n2550gat,
  II2414,n2633gat,II2417,n2551gat,II2420,n2552gat,II2425,n2553gat,II2428,
  n2554gat,II2433,n2555gat,II2439,n2545gat,n2619gat,n2504gat,n2660gat,
  n2655gat,n1528gat,n2293gat,n1523gat,n2219gat,n1592gat,n1529gat,n2666gat,
  n1704gat,n2422gat,n3013gat,n2290gat,n2081gat,n2218gat,n2285gat,n2359gat,
  n2358gat,n1414gat,n1415gat,n566gat,n1480gat,n2292gat,n1301gat,n1416gat,
  n1150gat,n873gat,n2011gat,n2306gat,n1478gat,n1481gat,n875gat,n1410gat,
  n2357gat,n876gat,n1347gat,n1160gat,n1484gat,n1084gat,n983gat,n1482gat,
  n2363gat,n1157gat,n1483gat,n985gat,n1530gat,n2364gat,n1307gat,n1308gat,
  n1085gat,n1479gat,n2291gat,n1348gat,n1349gat,n2217gat,n1591gat,n2223gat,
  n1437gat,n1438gat,n1832gat,n1765gat,n1878gat,n1442gat,n1831gat,n1444gat,
  n1378gat,n2975gat,n1322gat,n2974gat,n1439gat,n1486gat,n1370gat,n1426gat,
  n1369gat,n2966gat,n1366gat,n1365gat,n1374gat,n2979gat,n2162gat,n2220gat,
  n1450gat,n1423gat,n1427gat,n1608gat,n2082gat,n1449gat,n1494gat,n1590gat,
  n1248gat,n2954gat,n1418gat,n1417gat,n1306gat,n2964gat,n1353gat,n1419gat,
  n1247gat,n2958gat,n1355gat,n1422gat,n1300gat,n2963gat,n1487gat,n1485gat,
  n1164gat,n2953gat,n1356gat,n1354gat,n1436gat,n1435gat,n1106gat,n2949gat,
  n1425gat,n1421gat,n1105gat,n2934gat,n1424gat,n1420gat,n1309gat,n2959gat,
  II2672,n2142gat,n1788gat,II2684,n2060gat,n1786gat,II2696,n2138gat,n1839gat,
  n1897gat,n1884gat,n1848gat,n1783gat,n1548gat,II2721,n1719gat,n2137gat,
  n1633gat,n2059gat,n1785gat,II2731,n1849gat,n1784gat,n1716gat,II2736,
  n1635gat,n2401gat,n1989gat,n2392gat,n1918gat,II2771,n2439gat,n1986gat,
  n1866gat,n1865gat,II2785,n2406gat,n2216gat,n2345gat,n1988gat,n1735gat,
  n1861gat,n1387gat,n1694gat,II2813,n1780gat,n2019gat,n1549gat,II2832,
  n1551gat,II2837,n2346gat,n2152gat,n2405gat,n2351gat,II2843,n2402gat,
  n2212gat,II2847,n2393gat,n1991gat,n1665gat,n1666gat,n1517gat,n1578gat,
  II2873,n1495gat,n1604gat,II2885,n2090gat,n1550gat,II2890,n1552gat,n1738gat,
  II2915,n1739gat,n1925gat,n1920gat,n1917gat,n1921gat,n2141gat,n1787gat,
  II2926,n1859gat,n1922gat,n1798gat,II2935,n1743gat,n1923gat,n1864gat,
  n1690gat,II2953,n2178gat,n1661gat,n1660gat,n1572gat,n1576gat,n2438gat,
  n2283gat,n1520gat,n1582gat,n1580gat,n1577gat,n1990gat,n2988gat,II2978,
  n2189gat,II2989,n2134gat,II3000,n2261gat,n2128gat,n2129gat,n1695gat,II3016,
  n2181gat,II3056,n1311gat,n1707gat,n1659gat,n2987gat,n1515gat,n1521gat,
  n1736gat,n1737gat,n1658gat,n1724gat,n1732gat,n1662gat,n1663gat,n1656gat,
  n1655gat,n1670gat,n1667gat,n1569gat,n1570gat,n1568gat,n1575gat,n1727gat,
  n1728gat,n1797gat,n1801gat,n1730gat,n1731gat,n1561gat,n1571gat,n1668gat,
  n1734gat,n1742gat,n1671gat,n1669gat,n1652gat,n1657gat,n1648gat,n1729gat,
  n1790gat,n1726gat,n2004gat,n1929gat,n1869gat,II3143,n2591gat,n1584gat,
  n1714gat,II3149,n1718gat,II3163,n1507gat,n1396gat,n1401gat,II3168,n1393gat,
  n1409gat,n1476gat,II3174,n1898gat,n1838gat,II3179,II3191,n1677gat,n2000gat,
  n1412gat,n2001gat,n1999gat,II3211,n2663gat,n3018gat,n2448gat,n2662gat,
  n2444gat,II3235,n2238gat,n3019gat,n1310gat,n199gat,n87gat,n195gat,n184gat,
  n204gat,II3273,n2168gat,n2452gat,n1691gat,II3287,n3020gat,II3290,n3021gat,
  II3293,n3022gat,n1699gat,II3297,n3023gat,II3300,n3024gat,II3303,n3025gat,
  II3306,n3026gat,II3309,n3027gat,II3312,n3028gat,II3315,n3029gat,II3318,
  n3030gat,n2260gat,n2257gat,n2188gat,n2187gat,n3004gat,II3336,n2039gat,
  II3339,n1774gat,II3342,n1315gat,n2097gat,n1855gat,n2014gat,II3387,n2194gat,
  II3390,n3032gat,n2256gat,II3394,n3033gat,n2251gat,n2184gat,n3003gat,II3401,
  n2192gat,n2133gat,n2131gat,n2185gat,n2049gat,n3001gat,II3412,n2057gat,
  n2253gat,n2252gat,n2248gat,n3006gat,n2264gat,II3429,n2265gat,n2492gat,
  n2329gat,II3436,n1709gat,n1845gat,n1891gat,n1963gat,n1886gat,n1968gat,
  n1958gat,n1629gat,n1895gat,n1631gat,n1711gat,n2990gat,n2200gat,n2078gat,
  n2437gat,n2195gat,II3457,n2556gat,n1956gat,II3461,n3038gat,n1954gat,II3465,
  n3039gat,n1888gat,n2048gat,n2994gat,II3472,n2539gat,n1969gat,n1893gat,
  n1892gat,n2993gat,II3483,n2436gat,n2056gat,n2998gat,II3491,n2387gat,II3494,
  n3043gat,n1960gat,n1887gat,n1961gat,n2996gat,II3504,n2330gat,n2199gat,
  n2147gat,II3509,n3045gat,n2332gat,II3513,n3046gat,n2259gat,n2328gat,
  n3008gat,II3520,n2498gat,n2151gat,n2193gat,n2209gat,n3005gat,II3530,
  n2396gat,n2052gat,n2058gat,n2997gat,II3539,n2198gat,n2349gat,n2215gat,
  n2281gat,n3009gat,II3549,n2197gat,n2146gat,n3002gat,II3558,n2196gat,II3587,
  n2124gat,n2115gat,II3610,n1882gat,II3621,n1974gat,n1955gat,n1970gat,
  n1896gat,n1973gat,n2558gat,n2559gat,II3635,II3646,n2643gat,n2333gat,
  n2564gat,n2352gat,n2642gat,n2636gat,n2637gat,II3660,n88gat,n84gat,n375gat,
  n110gat,II3677,n155gat,n253gat,n1702gat,n150gat,II3691,n151gat,n243gat,
  n233gat,n154gat,n800gat,n2874gat,II3703,n2917gat,n235gat,n2878gat,II3713,
  n2892gat,n372gat,n212gat,n329gat,II3736,n387gat,n334gat,n1700gat,n386gat,
  II3742,n330gat,n1430gat,n1490gat,n452gat,n2885gat,II3754,n2900gat,n333gat,
  n2883gat,II3765,n2929gat,II3777,n462gat,n325gat,n457gat,n2884gat,n461gat,
  n458gat,n2902gat,II3801,n2925gat,n144gat,n247gat,II3808,n326gat,n878gat,
  n2879gat,II3817,n2916gat,n382gat,II3831,n383gat,n134gat,n2875gat,II3841,
  n2899gat,n254gat,n252gat,n2877gat,n468gat,II3867,n469gat,n381gat,n2893gat,
  II3876,n2926gat,n241gat,n140gat,II3882,n255gat,n802gat,n2882gat,II3891,
  n2924gat,n146gat,II3904,n147gat,n380gat,n2881gat,II3914,n2923gat,n69gat,
  n68gat,n1885gat,II3923,n2710gat,n2707gat,n16gat,n295gat,n357gat,n11gat,
  n12gat,n1889gat,II3935,n2704gat,n2700gat,n2051gat,II3941,n2684gat,n2680gat,
  n1350gat,II3945,n2696gat,II3948,n2692gat,II3951,n2683gat,II3954,n2679gat,
  II3957,n2449gat,n1754gat,II3962,n2830gat,n2827gat,n2512gat,n1544gat,
  n1769gat,n1683gat,n1756gat,n2167gat,n2013gat,II4000,n1791gat,n2691gat,
  n2695gat,n1518gat,n2699gat,n2703gat,n2159gat,n2478gat,II4014,n2744gat,
  n2740gat,n2158gat,n2186gat,II4020,n2800gat,n2797gat,n2288gat,II4024,
  n1513gat,n2537gat,n2538gat,n2442gat,n2483gat,n1334gat,II4055,n1747gat,
  II4067,n1674gat,n1403gat,n1402gat,II4081,n1806gat,n1634gat,n1338gat,II4105,
  n1455gat,II4108,n1339gat,n1505gat,n2980gat,II4117,n2758gat,n2755gat,
  n1546gat,II4122,n2752gat,n2748gat,n2012gat,n2016gat,n2002gat,n2008gat,
  II4129,n2858gat,n2857gat,II4135,n2766gat,II4138,n2765gat,n1684gat,n1759gat,
  II4145,II4157,n1524gat,n1862gat,n1863gat,n1919gat,n1860gat,n1460gat,II4185,
  n1595gat,n1454gat,n1469gat,n1468gat,n1519gat,II4194,n1461gat,n1477gat,
  n2984gat,n1594gat,II4212,n1587gat,n1681gat,II4217,II4222,n1761gat,n2751gat,
  n2747gat,II4227,n1760gat,n2743gat,n2739gat,n1978gat,II4233,n1721gat,
  n2808gat,II4236,n2804gat,n517gat,n518gat,n417gat,n418gat,n413gat,n411gat,
  n412gat,n522gat,n406gat,n516gat,n407gat,n355gat,n290gat,n525gat,n527gat,
  n356gat,n416gat,n415gat,n528gat,n521gat,n358gat,n532gat,n639gat,n523gat,
  n1111gat,n635gat,n524gat,n414gat,n1112gat,n630gat,n741gat,n629gat,n633gat,
  n634gat,n926gat,n632gat,n670gat,n636gat,n1123gat,n1007gat,n1006gat,II4309,
  n2941gat,n2814gat,II4312,n2811gat,n1002gat,n2946gat,II4329,n2950gat,
  n2813gat,II4332,n2810gat,n888gat,n2933gat,II4349,n2935gat,n2818gat,II4352,
  n2816gat,n898gat,n2940gat,II4369,n2937gat,n2817gat,II4372,n2815gat,
  n1179gat,n2947gat,II4389,n2956gat,n2824gat,II4392,n2821gat,n897gat,
  n2939gat,II4409,n2938gat,n2823gat,II4412,n2820gat,n894gat,n2932gat,II4429,
  n2936gat,n2829gat,II4432,n2826gat,n1180gat,n2948gat,II4449,n2955gat,
  n2828gat,II4452,n2825gat,n671gat,n628gat,n631gat,n976gat,II4475,n2951gat,
  n2807gat,II4478,n2803gat,n2127gat,II4482,n2682gat,II4485,n2678gat,n2046gat,
  II4489,n2681gat,II4492,n2677gat,n1708gat,II4496,n2688gat,II4499,n2686gat,
  n455gat,n291gat,n2237gat,II4506,n2764gat,n2763gat,n1782gat,II4512,n2762gat,
  n2760gat,n2325gat,II4518,n2761gat,n2759gat,n2245gat,II4524,n2757gat,
  n2754gat,n2244gat,II4530,n2756gat,n2753gat,n2243gat,II4536,n2750gat,
  n2746gat,n2246gat,II4542,n2749gat,n2745gat,n2384gat,II4548,n2742gat,
  n2738gat,n2385gat,II4554,n2741gat,n2737gat,n1286gat,II4558,n2687gat,
  n2685gat,n1328gat,n1381gat,n1384gat,II4566,n2694gat,n2690gat,n1382gat,
  n1451gat,n1453gat,II4573,n2693gat,n2689gat,n927gat,n925gat,n1452gat,II4580,
  n2702gat,n2698gat,n923gat,n921gat,n1890gat,II4587,n2701gat,n2697gat,
  n850gat,n739gat,n1841gat,II4594,n2709gat,n2706gat,n922gat,n848gat,n2047gat,
  II4601,n2708gat,n2705gat,n924gat,n849gat,n2050gat,II4608,n2799gat,n2796gat,
  n1118gat,n1032gat,n2054gat,II4615,n2798gat,n2795gat,II4620,n1745gat,
  n2806gat,II4623,n2802gat,II4626,n1870gat,n1086gat,II4630,n2805gat,II4633,
  n2801gat,n67gat,n85gat,n71gat,n180gat,n1840gat,II4642,n2812gat,n2809gat,
  n76gat,n82gat,n14gat,n186gat,n1842gat,II4651,n2822gat,n2819gat,II4654,
  II4657,II4660,II4663,II4666,II4669,II4672,II4675,II4678,II4681,II4684,
  II4687,II4690,II4693,II4696,II4699,II4702,II4705,II4708,II4711,II4714,
  II4717,II4720,II4723,II4726,II4729,II4732,II4735,II4738,II4741,II4744,
  II4747,II4750,II4753,II4756,II4759,II4762,II4765,II4768,II4771,II4774,
  II4777,II4780,II4783,II4786,II4789,II4792,II4795,II4798,n648gat,n442gat,
  n1214gat,n1215gat,n1216gat,n1217gat,n745gat,n638gat,n423gat,n362gat,
  n749gat,n750gat,n751gat,n752gat,n259gat,n260gat,n261gat,n262gat,n1014gat,
  n1015gat,n1016gat,n1017gat,n476gat,n477gat,n478gat,n479gat,n44gat,n45gat,
  n46gat,n47gat,n168gat,n169gat,n170gat,n171gat,n907gat,n908gat,n909gat,
  n910gat,n344gat,n345gat,n346gat,n347gat,n56gat,n57gat,n58gat,n59gat,
  n768gat,n655gat,n963gat,n868gat,n962gat,n959gat,n945gat,n946gat,n947gat,
  n948gat,n647gat,n441gat,n967gat,n792gat,n1229gat,n1230gat,n1231gat,
  n1232gat,n443gat,n439gat,n966gat,n790gat,n444gat,n440gat,n1051gat,n1052gat,
  n1053gat,n1054gat,n934gat,n935gat,n936gat,n937gat,n710gat,n711gat,n712gat,
  n713gat,n729gat,n730gat,n731gat,n732gat,n494gat,n495gat,n496gat,n497gat,
  n505gat,n506gat,n507gat,n508gat,II1277,n767gat,n653gat,n867gat,n771gat,
  n964gat,n961gat,n804gat,n805gat,n806gat,n807gat,n587gat,n588gat,n589gat,
  n590gat,n447gat,n445gat,n687gat,n688gat,n689gat,n690gat,n568gat,n569gat,
  n570gat,n571gat,II1515,II1584,n1692gat,II1723,II1733,n2428gat,n769gat,
  n1076gat,n766gat,n1185gat,n1186gat,n1187gat,n1188gat,n645gat,n646gat,
  n1383gat,n1327gat,n651gat,n652gat,n765gat,n1202gat,n1203gat,n1204gat,
  n1205gat,n1270gat,n1271gat,n1272gat,n1273gat,n763gat,n1287gat,n1285gat,
  n793gat,n556gat,n795gat,n656gat,n794gat,n773gat,n965gat,n960gat,n780gat,
  n781gat,n782gat,n783gat,n555gat,n450gat,n654gat,n557gat,n874gat,n132gat,
  n649gat,n449gat,n791gat,n650gat,n774gat,n764gat,n222gat,n223gat,n224gat,
  n225gat,n121gat,n122gat,n123gat,n124gat,n2460gat,n2423gat,n2569gat,
  n2570gat,n2571gat,n2572gat,n2410gat,n2411gat,n2412gat,n2413gat,n2580gat,
  n2581gat,n2567gat,n2499gat,n299gat,n207gat,n2647gat,n2648gat,n2602gat,
  n2603gat,n2604gat,n2605gat,n2546gat,n2547gat,n2548gat,n2549gat,n2614gat,
  n2615gat,n2461gat,n2421gat,n2930gat,n1153gat,n1151gat,n982gat,n877gat,
  n2957gat,n1159gat,n1158gat,n1156gat,n1155gat,n1443gat,n1325gat,n1321gat,
  n1320gat,n1368gat,n1258gat,n1373gat,n1372gat,n2978gat,n1441gat,n1440gat,
  n1371gat,n1367gat,n2982gat,n1504gat,n1502gat,n1250gat,n1103gat,n1304gat,
  n1249gat,n1246gat,n1161gat,n1291gat,n1245gat,n2973gat,n1352gat,n1351gat,
  n1303gat,n1302gat,n1163gat,n1102gat,n1101gat,n996gat,n1104gat,n887gat,
  n1305gat,n1162gat,n2977gat,n1360gat,n1359gat,n1358gat,n1357gat,II2720,
  II2735,II2812,n1703gat,n1778gat,n1609gat,II2831,II2889,II2925,II2934,
  n1733gat,n1581gat,n2079gat,n2073gat,n1574gat,n1573gat,n2992gat,n1723gat,
  n1647gat,n1646gat,n2986gat,n1650gat,n1649gat,n1563gat,n2991gat,n1654gat,
  n1653gat,n1644gat,II3148,II3178,n2981gat,n1413gat,n1408gat,n1407gat,
  n2258gat,n2255gat,n2132gat,n2130gat,n3007gat,n2250gat,n2249gat,n1710gat,
  n1630gat,n1894gat,n1847gat,n1846gat,n2055gat,n1967gat,n1959gat,n1957gat,
  n2211gat,n2210gat,n2053gat,n1964gat,n2350gat,n2282gat,n2213gat,n2150gat,
  n2149gat,n2995gat,n1962gat,n2999gat,n1972gat,n1971gat,n3011gat,n2331gat,
  n3015gat,n2566gat,n2565gat,n141gat,n38gat,n37gat,n1074gat,n872gat,n234gat,
  n137gat,n378gat,n377gat,n250gat,n249gat,n248gat,n869gat,n453gat,n448gat,
  n251gat,n244gat,n974gat,n973gat,n870gat,n246gat,n245gat,n460gat,n459gat,
  n975gat,n972gat,n969gat,n145gat,n143gat,n971gat,n970gat,n968gat,n142gat,
  n40gat,n39gat,n772gat,n451gat,n446gat,n139gat,n136gat,n391gat,n390gat,
  n1083gat,n1077gat,n242gat,n240gat,n871gat,n797gat,n324gat,n238gat,n237gat,
  n1082gat,n796gat,n1599gat,II3999,n1586gat,n1755gat,II4023,n1470gat,
  n1400gat,n1399gat,n1398gat,II4144,n1467gat,n1466gat,n2985gat,n1686gat,
  n1533gat,n1532gat,n1531gat,II4216,n2931gat,n1100gat,n994gat,n989gat,
  n880gat,n2943gat,n1012gat,n905gat,n1003gat,n902gat,n1099gat,n998gat,
  n995gat,n980gat,n2960gat,n1175gat,n1174gat,n1001gat,n999gat,n2969gat,
  n1323gat,n1264gat,n981gat,n890gat,n889gat,n886gat,n892gat,n891gat,n2942gat,
  n904gat,n903gat,n1152gat,n1092gat,n997gat,n993gat,n900gat,n895gat,n1094gat,
  n1093gat,n988gat,n984gat,n2965gat,n1267gat,n1257gat,n1178gat,n1116gat,
  n2961gat,n1375gat,n1324gat,n1091gat,n1088gat,n992gat,n987gat,n899gat,
  n896gat,n2967gat,n1262gat,n1260gat,n1098gat,n1090gat,n986gat,n885gat,
  n901gat,n893gat,n1097gat,n1089gat,n1087gat,n991gat,n2968gat,n1326gat,
  n1261gat,n1177gat,n1115gat,n2944gat,n977gat,n2945gat,n1096gat,n1095gat,
  n990gat,n979gat,n2962gat,n1176gat,n1173gat,n1004gat,n1000gat,n1029gat,
  n1028gat,n1031gat,n1030gat,n1011gat,n1181gat,n1010gat,n1005gat,n1182gat,
  n73gat,n70gat,n77gat,n13gat,n1935gat,n197gat,n22gat,n93gat,n2239gat,
  n2433gat,n2427gat,n2583gat,n2650gat,n2617gat,n1598gat,n1154gat,n1411gat,
  n1498gat,n1607gat,n1428gat,n1794gat,n1796gat,n1792gat,n1406gat,n2664gat,
  n1926gat,n1916gat,n1994gat,n1924gat,n1758gat,n200gat,n196gat,n2018gat,
  n89gat,n1471gat,n1472gat,n1600gat,n1397gat,n2005gat,n1818gat,n1510gat,
  n1459gat,n1458gat,n1602gat,n520gat,n519gat,n410gat,n354gat,n408gat,n526gat,
  n531gat,n530gat,n359gat,n420gat,n801gat,n879gat,n1255gat,n1009gat,n409gat,
  n292gat,n419gat,n1243gat,n1171gat,n1244gat,n1265gat,n1254gat,n1008gat,
  n1253gat,n1266gat,n1200gat,n1172gat,n1251gat,n1259gat,n1212gat,n1263gat,
  n978gat,n1199gat,n1252gat,n1757gat;

dff DFF_0(CK,n673gat,n2897gat);
dff DFF_1(CK,n398gat,n2782gat);
dff DFF_2(CK,n402gat,n2790gat);
dff DFF_3(CK,n919gat,n2670gat);
dff DFF_4(CK,n846gat,n2793gat);
dff DFF_5(CK,n394gat,n2782gat);
dff DFF_6(CK,n703gat,n2790gat);
dff DFF_7(CK,n722gat,n2670gat);
dff DFF_8(CK,n726gat,n2793gat);
dff DFF_9(CK,n2510gat,n748gat);
dff DFF_10(CK,n271gat,n2732gat);
dff DFF_11(CK,n160gat,n2776gat);
dff DFF_12(CK,n337gat,n2735gat);
dff DFF_13(CK,n842gat,n2673gat);
dff DFF_14(CK,n341gat,n2779gat);
dff DFF_15(CK,n2522gat,n43gat);
dff DFF_16(CK,n2472gat,n1620gat);
dff DFF_17(CK,n2319gat,n2470gat);
dff DFF_18(CK,n1821gat,n1827gat);
dff DFF_19(CK,n1825gat,n1827gat);
dff DFF_20(CK,n2029gat,n1816gat);
dff DFF_21(CK,n1829gat,n2027gat);
dff DFF_22(CK,n283gat,n2732gat);
dff DFF_23(CK,n165gat,n2776gat);
dff DFF_24(CK,n279gat,n2735gat);
dff DFF_25(CK,n1026gat,n2673gat);
dff DFF_26(CK,n275gat,n2779gat);
dff DFF_27(CK,n2476gat,n55gat);
dff DFF_28(CK,n1068gat,n2914gat);
dff DFF_29(CK,n957gat,n2928gat);
dff DFF_30(CK,n861gat,n2927gat);
dff DFF_31(CK,n1294gat,n2896gat);
dff DFF_32(CK,n1241gat,n2922gat);
dff DFF_33(CK,n1298gat,n2897gat);
dff DFF_34(CK,n865gat,n2894gat);
dff DFF_35(CK,n1080gat,n2921gat);
dff DFF_36(CK,n1148gat,n2895gat);
dff DFF_37(CK,n2468gat,n933gat);
dff DFF_38(CK,n618gat,n2790gat);
dff DFF_39(CK,n491gat,n2782gat);
dff DFF_40(CK,n622gat,n2793gat);
dff DFF_41(CK,n626gat,n2670gat);
dff DFF_42(CK,n834gat,n3064gat);
dff DFF_43(CK,n707gat,n3055gat);
dff DFF_44(CK,n838gat,n3063gat);
dff DFF_45(CK,n830gat,n3062gat);
dff DFF_46(CK,n614gat,n3056gat);
dff DFF_47(CK,n2526gat,n504gat);
dff DFF_48(CK,n680gat,n2913gat);
dff DFF_49(CK,n816gat,n2920gat);
dff DFF_50(CK,n580gat,n2905gat);
dff DFF_51(CK,n824gat,n3057gat);
dff DFF_52(CK,n820gat,n3059gat);
dff DFF_53(CK,n883gat,n3058gat);
dff DFF_54(CK,n584gat,n2898gat);
dff DFF_55(CK,n684gat,n3060gat);
dff DFF_56(CK,n699gat,n3061gat);
dff DFF_57(CK,n2464gat,n567gat);
dff DFF_58(CK,n2399gat,n3048gat);
dff DFF_59(CK,n2343gat,n3049gat);
dff DFF_60(CK,n2203gat,n3051gat);
dff DFF_61(CK,n2562gat,n3047gat);
dff DFF_62(CK,n2207gat,n3050gat);
dff DFF_63(CK,n2626gat,n3040gat);
dff DFF_64(CK,n2490gat,n3044gat);
dff DFF_65(CK,n2622gat,n3042gat);
dff DFF_66(CK,n2630gat,n3037gat);
dff DFF_67(CK,n2543gat,n3041gat);
dff DFF_68(CK,n2102gat,n1606gat);
dff DFF_69(CK,n1880gat,n3052gat);
dff DFF_70(CK,n1763gat,n1610gat);
dff DFF_71(CK,n2155gat,n1858gat);
dff DFF_72(CK,n1035gat,n2918gat);
dff DFF_73(CK,n1121gat,n2952gat);
dff DFF_74(CK,n1072gat,n2919gat);
dff DFF_75(CK,n1282gat,n2910gat);
dff DFF_76(CK,n1226gat,n2907gat);
dff DFF_77(CK,n931gat,n2911gat);
dff DFF_78(CK,n1135gat,n2912gat);
dff DFF_79(CK,n1045gat,n2909gat);
dff DFF_80(CK,n1197gat,n2908gat);
dff DFF_81(CK,n2518gat,n2971gat);
dff DFF_82(CK,n667gat,n2904gat);
dff DFF_83(CK,n659gat,n2891gat);
dff DFF_84(CK,n553gat,n2903gat);
dff DFF_85(CK,n777gat,n2915gat);
dff DFF_86(CK,n561gat,n2901gat);
dff DFF_87(CK,n366gat,n2890gat);
dff DFF_88(CK,n322gat,n2888gat);
dff DFF_89(CK,n318gat,n2887gat);
dff DFF_90(CK,n314gat,n2886gat);
dff DFF_91(CK,n2599gat,n3010gat);
dff DFF_92(CK,n2588gat,n3016gat);
dff DFF_93(CK,n2640gat,n3054gat);
dff DFF_94(CK,n2658gat,n2579gat);
dff DFF_95(CK,n2495gat,n3036gat);
dff DFF_96(CK,n2390gat,n3034gat);
dff DFF_97(CK,n2270gat,n3031gat);
dff DFF_98(CK,n2339gat,n3035gat);
dff DFF_99(CK,n2502gat,n2646gat);
dff DFF_100(CK,n2634gat,n3053gat);
dff DFF_101(CK,n2506gat,n2613gat);
dff DFF_102(CK,n1834gat,n1625gat);
dff DFF_103(CK,n1767gat,n1626gat);
dff DFF_104(CK,n2084gat,n1603gat);
dff DFF_105(CK,n2143gat,n2541gat);
dff DFF_106(CK,n2061gat,n2557gat);
dff DFF_107(CK,n2139gat,n2487gat);
dff DFF_108(CK,n1899gat,n2532gat);
dff DFF_109(CK,n1850gat,n2628gat);
dff DFF_110(CK,n2403gat,n2397gat);
dff DFF_111(CK,n2394gat,n2341gat);
dff DFF_112(CK,n2440gat,n2560gat);
dff DFF_113(CK,n2407gat,n2205gat);
dff DFF_114(CK,n2347gat,n2201gat);
dff DFF_115(CK,n1389gat,n1793gat);
dff DFF_116(CK,n2021gat,n1781gat);
dff DFF_117(CK,n1394gat,n1516gat);
dff DFF_118(CK,n1496gat,n1392gat);
dff DFF_119(CK,n2091gat,n1685gat);
dff DFF_120(CK,n1332gat,n1565gat);
dff DFF_121(CK,n1740gat,n1330gat);
dff DFF_122(CK,n2179gat,n1945gat);
dff DFF_123(CK,n2190gat,n2268gat);
dff DFF_124(CK,n2135gat,n2337gat);
dff DFF_125(CK,n2262gat,n2388gat);
dff DFF_126(CK,n2182gat,n1836gat);
dff DFF_127(CK,n1433gat,n2983gat);
dff DFF_128(CK,n1316gat,n1431gat);
dff DFF_129(CK,n1363gat,n1314gat);
dff DFF_130(CK,n1312gat,n1361gat);
dff DFF_131(CK,n1775gat,n1696gat);
dff DFF_132(CK,n1871gat,n2009gat);
dff DFF_133(CK,n2592gat,n1773gat);
dff DFF_134(CK,n1508gat,n1636gat);
dff DFF_135(CK,n1678gat,n1712gat);
dff DFF_136(CK,n2309gat,n3000gat);
dff DFF_137(CK,n2450gat,n2307gat);
dff DFF_138(CK,n2446gat,n2661gat);
dff DFF_139(CK,n2095gat,n827gat);
dff DFF_140(CK,n2176gat,n2093gat);
dff DFF_141(CK,n2169gat,n2174gat);
dff DFF_142(CK,n2454gat,n2163gat);
dff DFF_143(CK,n2040gat,n1777gat);
dff DFF_144(CK,n2044gat,n2015gat);
dff DFF_145(CK,n2037gat,n2042gat);
dff DFF_146(CK,n2025gat,n2017gat);
dff DFF_147(CK,n2099gat,n2023gat);
dff DFF_148(CK,n2266gat,n2493gat);
dff DFF_149(CK,n2033gat,n2035gat);
dff DFF_150(CK,n2110gat,n2031gat);
dff DFF_151(CK,n2125gat,n2108gat);
dff DFF_152(CK,n2121gat,n2123gat);
dff DFF_153(CK,n2117gat,n2119gat);
dff DFF_154(CK,n1975gat,n2632gat);
dff DFF_155(CK,n2644gat,n2638gat);
dff DFF_156(CK,n156gat,n612gat);
dff DFF_157(CK,n152gat,n705gat);
dff DFF_158(CK,n331gat,n822gat);
dff DFF_159(CK,n388gat,n881gat);
dff DFF_160(CK,n463gat,n818gat);
dff DFF_161(CK,n327gat,n682gat);
dff DFF_162(CK,n384gat,n697gat);
dff DFF_163(CK,n256gat,n836gat);
dff DFF_164(CK,n470gat,n828gat);
dff DFF_165(CK,n148gat,n832gat);
dff DFF_166(CK,n2458gat,n2590gat);
dff DFF_167(CK,n2514gat,n2456gat);
dff DFF_168(CK,n1771gat,n1613gat);
dff DFF_169(CK,n1336gat,n1391gat);
dff DFF_170(CK,n1748gat,n1927gat);
dff DFF_171(CK,n1675gat,n1713gat);
dff DFF_172(CK,n1807gat,n1717gat);
dff DFF_173(CK,n1340gat,n1567gat);
dff DFF_174(CK,n1456gat,n1564gat);
dff DFF_175(CK,n1525gat,n1632gat);
dff DFF_176(CK,n1462gat,n1915gat);
dff DFF_177(CK,n1596gat,n1800gat);
dff DFF_178(CK,n1588gat,n1593gat);
not NOT_0(II1,n3088gat);
not NOT_1(n2717gat,II1);
not NOT_2(n2715gat,n2717gat);
not NOT_3(II5,n3087gat);
not NOT_4(n2725gat,II5);
not NOT_5(n2723gat,n2725gat);
not NOT_6(n296gat,n421gat);
not NOT_7(II11,n3093gat);
not NOT_8(n2768gat,II11);
not NOT_9(II14,n2768gat);
not NOT_10(n2767gat,II14);
not NOT_11(n373gat,n2767gat);
not NOT_12(II18,n3072gat);
not NOT_13(n2671gat,II18);
not NOT_14(n2669gat,n2671gat);
not NOT_15(II23,n3081gat);
not NOT_16(n2845gat,II23);
not NOT_17(n2844gat,n2845gat);
not NOT_18(II27,n3095gat);
not NOT_19(n2668gat,II27);
not NOT_20(II30,n2668gat);
not NOT_21(n2667gat,II30);
not NOT_22(n856gat,n2667gat);
not NOT_23(II44,n673gat);
not NOT_24(n672gat,II44);
not NOT_25(II47,n3069gat);
not NOT_26(n2783gat,II47);
not NOT_27(II50,n2783gat);
not NOT_28(n2782gat,II50);
not NOT_29(n396gat,n398gat);
not NOT_30(II62,n3070gat);
not NOT_31(n2791gat,II62);
not NOT_32(II65,n2791gat);
not NOT_33(n2790gat,II65);
not NOT_34(II76,n402gat);
not NOT_35(n401gat,II76);
not NOT_36(n1645gat,n1499gat);
not NOT_37(II81,n2671gat);
not NOT_38(n2670gat,II81);
not NOT_39(II92,n919gat);
not NOT_40(n918gat,II92);
not NOT_41(n1553gat,n1616gat);
not NOT_42(II97,n3071gat);
not NOT_43(n2794gat,II97);
not NOT_44(II100,n2794gat);
not NOT_45(n2793gat,II100);
not NOT_46(II111,n846gat);
not NOT_47(n845gat,II111);
not NOT_48(n1559gat,n1614gat);
not NOT_49(n1643gat,n1641gat);
not NOT_50(n1651gat,n1642gat);
not NOT_51(n1562gat,n1556gat);
not NOT_52(n1560gat,n1557gat);
not NOT_53(n1640gat,n1639gat);
not NOT_54(n1566gat,n1605gat);
not NOT_55(n1554gat,n1555gat);
not NOT_56(n1722gat,n1558gat);
not NOT_57(n392gat,n394gat);
not NOT_58(II149,n703gat);
not NOT_59(n702gat,II149);
not NOT_60(n1319gat,n1256gat);
not NOT_61(n720gat,n722gat);
not NOT_62(II171,n726gat);
not NOT_63(n725gat,II171);
not NOT_64(n1447gat,n1117gat);
not NOT_65(n1627gat,n1618gat);
not NOT_66(II178,n722gat);
not NOT_67(n721gat,II178);
not NOT_68(n1380gat,n1114gat);
not NOT_69(n1628gat,n1621gat);
not NOT_70(n701gat,n703gat);
not NOT_71(n1446gat,n1318gat);
not NOT_72(n1705gat,n1619gat);
not NOT_73(n1706gat,n1622gat);
not NOT_74(II192,n3083gat);
not NOT_75(n2856gat,II192);
not NOT_76(n2854gat,n2856gat);
not NOT_77(II196,n2854gat);
not NOT_78(n1218gat,II196);
not NOT_79(II199,n3085gat);
not NOT_80(n2861gat,II199);
not NOT_81(n2859gat,n2861gat);
not NOT_82(II203,n2859gat);
not NOT_83(n1219gat,II203);
not NOT_84(II206,n3084gat);
not NOT_85(n2864gat,II206);
not NOT_86(n2862gat,n2864gat);
not NOT_87(II210,n2862gat);
not NOT_88(n1220gat,II210);
not NOT_89(II214,n2861gat);
not NOT_90(n2860gat,II214);
not NOT_91(II217,n2860gat);
not NOT_92(n1221gat,II217);
not NOT_93(II220,n2864gat);
not NOT_94(n2863gat,II220);
not NOT_95(II223,n2863gat);
not NOT_96(n1222gat,II223);
not NOT_97(II227,n2856gat);
not NOT_98(n2855gat,II227);
not NOT_99(II230,n2855gat);
not NOT_100(n1223gat,II230);
not NOT_101(n640gat,n1213gat);
not NOT_102(II237,n640gat);
not NOT_103(n753gat,II237);
not NOT_104(II240,n2717gat);
not NOT_105(n2716gat,II240);
not NOT_106(II243,n3089gat);
not NOT_107(n2869gat,II243);
not NOT_108(n2867gat,n2869gat);
not NOT_109(II248,n2869gat);
not NOT_110(n2868gat,II248);
not NOT_111(II253,n2906gat);
not NOT_112(n754gat,II253);
not NOT_113(II256,n2725gat);
not NOT_114(n2724gat,II256);
not NOT_115(II259,n3086gat);
not NOT_116(n2728gat,II259);
not NOT_117(n2726gat,n2728gat);
not NOT_118(II264,n2728gat);
not NOT_119(n2727gat,II264);
not NOT_120(n422gat,n2889gat);
not NOT_121(II270,n422gat);
not NOT_122(n755gat,II270);
not NOT_123(n747gat,n2906gat);
not NOT_124(II275,n747gat);
not NOT_125(n756gat,II275);
not NOT_126(II278,n2889gat);
not NOT_127(n757gat,II278);
not NOT_128(II282,n1213gat);
not NOT_129(n758gat,II282);
not NOT_130(n2508gat,n2510gat);
not NOT_131(II297,n3065gat);
not NOT_132(n2733gat,II297);
not NOT_133(II300,n2733gat);
not NOT_134(n2732gat,II300);
not NOT_135(II311,n271gat);
not NOT_136(n270gat,II311);
not NOT_137(II314,n270gat);
not NOT_138(n263gat,II314);
not NOT_139(II317,n3067gat);
not NOT_140(n2777gat,II317);
not NOT_141(II320,n2777gat);
not NOT_142(n2776gat,II320);
not NOT_143(II331,n160gat);
not NOT_144(n159gat,II331);
not NOT_145(II334,n159gat);
not NOT_146(n264gat,II334);
not NOT_147(II337,n3066gat);
not NOT_148(n2736gat,II337);
not NOT_149(II340,n2736gat);
not NOT_150(n2735gat,II340);
not NOT_151(II351,n337gat);
not NOT_152(n336gat,II351);
not NOT_153(II354,n336gat);
not NOT_154(n265gat,II354);
not NOT_155(n158gat,n160gat);
not NOT_156(II359,n158gat);
not NOT_157(n266gat,II359);
not NOT_158(n335gat,n337gat);
not NOT_159(II363,n335gat);
not NOT_160(n267gat,II363);
not NOT_161(n269gat,n271gat);
not NOT_162(II368,n269gat);
not NOT_163(n268gat,II368);
not NOT_164(n41gat,n258gat);
not NOT_165(II375,n41gat);
not NOT_166(n48gat,II375);
not NOT_167(II378,n725gat);
not NOT_168(n1018gat,II378);
not NOT_169(II381,n3073gat);
not NOT_170(n2674gat,II381);
not NOT_171(II384,n2674gat);
not NOT_172(n2673gat,II384);
not NOT_173(II395,n842gat);
not NOT_174(n841gat,II395);
not NOT_175(II398,n841gat);
not NOT_176(n1019gat,II398);
not NOT_177(II401,n721gat);
not NOT_178(n1020gat,II401);
not NOT_179(n840gat,n842gat);
not NOT_180(II406,n840gat);
not NOT_181(n1021gat,II406);
not NOT_182(II409,n720gat);
not NOT_183(n1022gat,II409);
not NOT_184(n724gat,n726gat);
not NOT_185(II414,n724gat);
not NOT_186(n1023gat,II414);
not NOT_187(II420,n1013gat);
not NOT_188(n49gat,II420);
not NOT_189(II423,n3068gat);
not NOT_190(n2780gat,II423);
not NOT_191(II426,n2780gat);
not NOT_192(n2779gat,II426);
not NOT_193(II437,n341gat);
not NOT_194(n340gat,II437);
not NOT_195(II440,n340gat);
not NOT_196(n480gat,II440);
not NOT_197(II443,n702gat);
not NOT_198(n481gat,II443);
not NOT_199(II446,n394gat);
not NOT_200(n393gat,II446);
not NOT_201(II449,n393gat);
not NOT_202(n482gat,II449);
not NOT_203(II453,n701gat);
not NOT_204(n483gat,II453);
not NOT_205(II456,n392gat);
not NOT_206(n484gat,II456);
not NOT_207(n339gat,n341gat);
not NOT_208(II461,n339gat);
not NOT_209(n485gat,II461);
not NOT_210(n42gat,n475gat);
not NOT_211(II468,n42gat);
not NOT_212(n50gat,II468);
not NOT_213(n162gat,n1013gat);
not NOT_214(II473,n162gat);
not NOT_215(n51gat,II473);
not NOT_216(II476,n475gat);
not NOT_217(n52gat,II476);
not NOT_218(II480,n258gat);
not NOT_219(n53gat,II480);
not NOT_220(n2520gat,n2522gat);
not NOT_221(n1448gat,n1376gat);
not NOT_222(n1701gat,n1617gat);
not NOT_223(n1379gat,n1377gat);
not NOT_224(n1615gat,n1624gat);
not NOT_225(n1500gat,n1113gat);
not NOT_226(n1503gat,n1501gat);
not NOT_227(n1779gat,n1623gat);
not NOT_228(II509,n3099gat);
not NOT_229(n2730gat,II509);
not NOT_230(II512,n2730gat);
not NOT_231(n2729gat,II512);
not NOT_232(n2470gat,n2472gat);
not NOT_233(n2317gat,n2319gat);
not NOT_234(n1819gat,n1821gat);
not NOT_235(n1823gat,n1825gat);
not NOT_236(n1816gat,n1817gat);
not NOT_237(n2027gat,n2029gat);
not NOT_238(II572,n1829gat);
not NOT_239(n1828gat,II572);
not NOT_240(II576,n3100gat);
not NOT_241(n2851gat,II576);
not NOT_242(II579,n2851gat);
not NOT_243(n2850gat,II579);
not NOT_244(II583,n2786gat);
not NOT_245(n2785gat,II583);
not NOT_246(n92gat,n2785gat);
not NOT_247(n637gat,n529gat);
not NOT_248(n293gat,n361gat);
not NOT_249(II591,n3094gat);
not NOT_250(n2722gat,II591);
not NOT_251(II594,n2722gat);
not NOT_252(n2721gat,II594);
not NOT_253(n297gat,n2721gat);
not NOT_254(II606,n283gat);
not NOT_255(n282gat,II606);
not NOT_256(II609,n282gat);
not NOT_257(n172gat,II609);
not NOT_258(II620,n165gat);
not NOT_259(n164gat,II620);
not NOT_260(II623,n164gat);
not NOT_261(n173gat,II623);
not NOT_262(II634,n279gat);
not NOT_263(n278gat,II634);
not NOT_264(II637,n278gat);
not NOT_265(n174gat,II637);
not NOT_266(n163gat,n165gat);
not NOT_267(II642,n163gat);
not NOT_268(n175gat,II642);
not NOT_269(n277gat,n279gat);
not NOT_270(II646,n277gat);
not NOT_271(n176gat,II646);
not NOT_272(n281gat,n283gat);
not NOT_273(II651,n281gat);
not NOT_274(n177gat,II651);
not NOT_275(n54gat,n167gat);
not NOT_276(II658,n54gat);
not NOT_277(n60gat,II658);
not NOT_278(II661,n845gat);
not NOT_279(n911gat,II661);
not NOT_280(II672,n1026gat);
not NOT_281(n1025gat,II672);
not NOT_282(II675,n1025gat);
not NOT_283(n912gat,II675);
not NOT_284(II678,n918gat);
not NOT_285(n913gat,II678);
not NOT_286(n1024gat,n1026gat);
not NOT_287(II683,n1024gat);
not NOT_288(n914gat,II683);
not NOT_289(n917gat,n919gat);
not NOT_290(II687,n917gat);
not NOT_291(n915gat,II687);
not NOT_292(n844gat,n846gat);
not NOT_293(II692,n844gat);
not NOT_294(n916gat,II692);
not NOT_295(II698,n906gat);
not NOT_296(n61gat,II698);
not NOT_297(II709,n275gat);
not NOT_298(n274gat,II709);
not NOT_299(II712,n274gat);
not NOT_300(n348gat,II712);
not NOT_301(II715,n401gat);
not NOT_302(n349gat,II715);
not NOT_303(II718,n398gat);
not NOT_304(n397gat,II718);
not NOT_305(II721,n397gat);
not NOT_306(n350gat,II721);
not NOT_307(n400gat,n402gat);
not NOT_308(II726,n400gat);
not NOT_309(n351gat,II726);
not NOT_310(II729,n396gat);
not NOT_311(n352gat,II729);
not NOT_312(n273gat,n275gat);
not NOT_313(II734,n273gat);
not NOT_314(n353gat,II734);
not NOT_315(n178gat,n343gat);
not NOT_316(II741,n178gat);
not NOT_317(n62gat,II741);
not NOT_318(n66gat,n906gat);
not NOT_319(II746,n66gat);
not NOT_320(n63gat,II746);
not NOT_321(II749,n343gat);
not NOT_322(n64gat,II749);
not NOT_323(II753,n167gat);
not NOT_324(n65gat,II753);
not NOT_325(n2474gat,n2476gat);
not NOT_326(II768,n3090gat);
not NOT_327(n2832gat,II768);
not NOT_328(II771,n2832gat);
not NOT_329(n2831gat,II771);
not NOT_330(n2731gat,n2733gat);
not NOT_331(II776,n3074gat);
not NOT_332(n2719gat,II776);
not NOT_333(n2718gat,n2719gat);
not NOT_334(II790,n1068gat);
not NOT_335(n1067gat,II790);
not NOT_336(II793,n1067gat);
not NOT_337(n949gat,II793);
not NOT_338(II796,n3076gat);
not NOT_339(n2839gat,II796);
not NOT_340(n2838gat,n2839gat);
not NOT_341(n2775gat,n2777gat);
not NOT_342(II812,n957gat);
not NOT_343(n956gat,II812);
not NOT_344(II815,n956gat);
not NOT_345(n950gat,II815);
not NOT_346(II818,n3075gat);
not NOT_347(n2712gat,II818);
not NOT_348(n2711gat,n2712gat);
not NOT_349(n2734gat,n2736gat);
not NOT_350(II834,n861gat);
not NOT_351(n860gat,II834);
not NOT_352(II837,n860gat);
not NOT_353(n951gat,II837);
not NOT_354(n955gat,n957gat);
not NOT_355(II842,n955gat);
not NOT_356(n952gat,II842);
not NOT_357(n859gat,n861gat);
not NOT_358(II846,n859gat);
not NOT_359(n953gat,II846);
not NOT_360(n1066gat,n1068gat);
not NOT_361(II851,n1066gat);
not NOT_362(n954gat,II851);
not NOT_363(n857gat,n944gat);
not NOT_364(II858,n857gat);
not NOT_365(n938gat,II858);
not NOT_366(n2792gat,n2794gat);
not NOT_367(II863,n3080gat);
not NOT_368(n2847gat,II863);
not NOT_369(n2846gat,n2847gat);
not NOT_370(II877,n1294gat);
not NOT_371(n1293gat,II877);
not NOT_372(II880,n1293gat);
not NOT_373(n1233gat,II880);
not NOT_374(n2672gat,n2674gat);
not NOT_375(II885,n3082gat);
not NOT_376(n2853gat,II885);
not NOT_377(n2852gat,n2853gat);
not NOT_378(II899,n1241gat);
not NOT_379(n1240gat,II899);
not NOT_380(II902,n1240gat);
not NOT_381(n1234gat,II902);
not NOT_382(II913,n1298gat);
not NOT_383(n1297gat,II913);
not NOT_384(II916,n1297gat);
not NOT_385(n1235gat,II916);
not NOT_386(n1239gat,n1241gat);
not NOT_387(II921,n1239gat);
not NOT_388(n1236gat,II921);
not NOT_389(n1296gat,n1298gat);
not NOT_390(II925,n1296gat);
not NOT_391(n1237gat,II925);
not NOT_392(n1292gat,n1294gat);
not NOT_393(II930,n1292gat);
not NOT_394(n1238gat,II930);
not NOT_395(II936,n1228gat);
not NOT_396(n939gat,II936);
not NOT_397(n2778gat,n2780gat);
not NOT_398(II941,n3077gat);
not NOT_399(n2837gat,II941);
not NOT_400(n2836gat,n2837gat);
not NOT_401(II955,n865gat);
not NOT_402(n864gat,II955);
not NOT_403(II958,n864gat);
not NOT_404(n1055gat,II958);
not NOT_405(n2789gat,n2791gat);
not NOT_406(II963,n3079gat);
not NOT_407(n2841gat,II963);
not NOT_408(n2840gat,n2841gat);
not NOT_409(II977,n1080gat);
not NOT_410(n1079gat,II977);
not NOT_411(II980,n1079gat);
not NOT_412(n1056gat,II980);
not NOT_413(n2781gat,n2783gat);
not NOT_414(II985,n3078gat);
not NOT_415(n2843gat,II985);
not NOT_416(n2842gat,n2843gat);
not NOT_417(II999,n1148gat);
not NOT_418(n1147gat,II999);
not NOT_419(II1002,n1147gat);
not NOT_420(n1057gat,II1002);
not NOT_421(n1078gat,n1080gat);
not NOT_422(II1007,n1078gat);
not NOT_423(n1058gat,II1007);
not NOT_424(n1146gat,n1148gat);
not NOT_425(II1011,n1146gat);
not NOT_426(n1059gat,II1011);
not NOT_427(n863gat,n865gat);
not NOT_428(II1016,n863gat);
not NOT_429(n1060gat,II1016);
not NOT_430(n928gat,n1050gat);
not NOT_431(II1023,n928gat);
not NOT_432(n940gat,II1023);
not NOT_433(n858gat,n1228gat);
not NOT_434(II1028,n858gat);
not NOT_435(n941gat,II1028);
not NOT_436(II1031,n1050gat);
not NOT_437(n942gat,II1031);
not NOT_438(II1035,n944gat);
not NOT_439(n943gat,II1035);
not NOT_440(n2466gat,n2468gat);
not NOT_441(n2720gat,n2722gat);
not NOT_442(n740gat,n2667gat);
not NOT_443(n2784gat,n2786gat);
not NOT_444(n743gat,n746gat);
not NOT_445(n294gat,n360gat);
not NOT_446(n374gat,n2767gat);
not NOT_447(n616gat,n618gat);
not NOT_448(II1067,n616gat);
not NOT_449(n501gat,II1067);
not NOT_450(n489gat,n491gat);
not NOT_451(II1079,n489gat);
not NOT_452(n502gat,II1079);
not NOT_453(II1082,n618gat);
not NOT_454(n617gat,II1082);
not NOT_455(II1085,n617gat);
not NOT_456(n499gat,II1085);
not NOT_457(II1088,n491gat);
not NOT_458(n490gat,II1088);
not NOT_459(II1091,n490gat);
not NOT_460(n500gat,II1091);
not NOT_461(n620gat,n622gat);
not NOT_462(II1103,n620gat);
not NOT_463(n738gat,II1103);
not NOT_464(n624gat,n626gat);
not NOT_465(II1115,n624gat);
not NOT_466(n737gat,II1115);
not NOT_467(II1118,n622gat);
not NOT_468(n621gat,II1118);
not NOT_469(II1121,n621gat);
not NOT_470(n733gat,II1121);
not NOT_471(II1124,n626gat);
not NOT_472(n625gat,II1124);
not NOT_473(II1127,n625gat);
not NOT_474(n735gat,II1127);
not NOT_475(II1138,n834gat);
not NOT_476(n833gat,II1138);
not NOT_477(II1141,n833gat);
not NOT_478(n714gat,II1141);
not NOT_479(II1152,n707gat);
not NOT_480(n706gat,II1152);
not NOT_481(II1155,n706gat);
not NOT_482(n715gat,II1155);
not NOT_483(II1166,n838gat);
not NOT_484(n837gat,II1166);
not NOT_485(II1169,n837gat);
not NOT_486(n716gat,II1169);
not NOT_487(n705gat,n707gat);
not NOT_488(II1174,n705gat);
not NOT_489(n717gat,II1174);
not NOT_490(n836gat,n838gat);
not NOT_491(II1178,n836gat);
not NOT_492(n718gat,II1178);
not NOT_493(n832gat,n834gat);
not NOT_494(II1183,n832gat);
not NOT_495(n719gat,II1183);
not NOT_496(n515gat,n709gat);
not NOT_497(II1190,n515gat);
not NOT_498(n509gat,II1190);
not NOT_499(II1201,n830gat);
not NOT_500(n829gat,II1201);
not NOT_501(II1204,n829gat);
not NOT_502(n734gat,II1204);
not NOT_503(n828gat,n830gat);
not NOT_504(II1209,n828gat);
not NOT_505(n736gat,II1209);
not NOT_506(II1216,n728gat);
not NOT_507(n510gat,II1216);
not NOT_508(II1227,n614gat);
not NOT_509(n613gat,II1227);
not NOT_510(II1230,n613gat);
not NOT_511(n498gat,II1230);
not NOT_512(n612gat,n614gat);
not NOT_513(II1236,n612gat);
not NOT_514(n503gat,II1236);
not NOT_515(n404gat,n493gat);
not NOT_516(II1243,n404gat);
not NOT_517(n511gat,II1243);
not NOT_518(n405gat,n728gat);
not NOT_519(II1248,n405gat);
not NOT_520(n512gat,II1248);
not NOT_521(II1251,n493gat);
not NOT_522(n513gat,II1251);
not NOT_523(II1255,n709gat);
not NOT_524(n514gat,II1255);
not NOT_525(n2524gat,n2526gat);
not NOT_526(n17gat,n564gat);
not NOT_527(n79gat,n86gat);
not NOT_528(n219gat,n78gat);
not NOT_529(n563gat,II1278);
not NOT_530(n289gat,n563gat);
not NOT_531(n179gat,n287gat);
not NOT_532(n188gat,n288gat);
not NOT_533(n72gat,n181gat);
not NOT_534(n111gat,n182gat);
not NOT_535(II1302,n680gat);
not NOT_536(n679gat,II1302);
not NOT_537(II1305,n679gat);
not NOT_538(n808gat,II1305);
not NOT_539(II1319,n816gat);
not NOT_540(n815gat,II1319);
not NOT_541(II1322,n815gat);
not NOT_542(n809gat,II1322);
not NOT_543(II1336,n580gat);
not NOT_544(n579gat,II1336);
not NOT_545(II1339,n579gat);
not NOT_546(n810gat,II1339);
not NOT_547(n814gat,n816gat);
not NOT_548(II1344,n814gat);
not NOT_549(n811gat,II1344);
not NOT_550(n578gat,n580gat);
not NOT_551(II1348,n578gat);
not NOT_552(n812gat,II1348);
not NOT_553(n678gat,n680gat);
not NOT_554(II1353,n678gat);
not NOT_555(n813gat,II1353);
not NOT_556(n677gat,n803gat);
not NOT_557(II1360,n677gat);
not NOT_558(n572gat,II1360);
not NOT_559(II1371,n824gat);
not NOT_560(n823gat,II1371);
not NOT_561(II1374,n823gat);
not NOT_562(n591gat,II1374);
not NOT_563(II1385,n820gat);
not NOT_564(n819gat,II1385);
not NOT_565(II1388,n819gat);
not NOT_566(n592gat,II1388);
not NOT_567(II1399,n883gat);
not NOT_568(n882gat,II1399);
not NOT_569(II1402,n882gat);
not NOT_570(n593gat,II1402);
not NOT_571(n818gat,n820gat);
not NOT_572(II1407,n818gat);
not NOT_573(n594gat,II1407);
not NOT_574(n881gat,n883gat);
not NOT_575(II1411,n881gat);
not NOT_576(n595gat,II1411);
not NOT_577(n822gat,n824gat);
not NOT_578(II1416,n822gat);
not NOT_579(n596gat,II1416);
not NOT_580(II1422,n586gat);
not NOT_581(n573gat,II1422);
not NOT_582(II1436,n584gat);
not NOT_583(n583gat,II1436);
not NOT_584(II1439,n583gat);
not NOT_585(n691gat,II1439);
not NOT_586(II1450,n684gat);
not NOT_587(n683gat,II1450);
not NOT_588(II1453,n683gat);
not NOT_589(n692gat,II1453);
not NOT_590(II1464,n699gat);
not NOT_591(n698gat,II1464);
not NOT_592(II1467,n698gat);
not NOT_593(n693gat,II1467);
not NOT_594(n682gat,n684gat);
not NOT_595(II1472,n682gat);
not NOT_596(n694gat,II1472);
not NOT_597(n697gat,n699gat);
not NOT_598(II1476,n697gat);
not NOT_599(n695gat,II1476);
not NOT_600(n582gat,n584gat);
not NOT_601(II1481,n582gat);
not NOT_602(n696gat,II1481);
not NOT_603(n456gat,n686gat);
not NOT_604(II1488,n456gat);
not NOT_605(n574gat,II1488);
not NOT_606(n565gat,n586gat);
not NOT_607(II1493,n565gat);
not NOT_608(n575gat,II1493);
not NOT_609(II1496,n686gat);
not NOT_610(n576gat,II1496);
not NOT_611(II1500,n803gat);
not NOT_612(n577gat,II1500);
not NOT_613(n2462gat,n2464gat);
not NOT_614(n2665gat,II1516);
not NOT_615(n2596gat,n2665gat);
not NOT_616(n189gat,n286gat);
not NOT_617(n194gat,n187gat);
not NOT_618(n21gat,n15gat);
not NOT_619(II1538,n2399gat);
not NOT_620(n2398gat,II1538);
not NOT_621(n2353gat,n2398gat);
not NOT_622(II1550,n2343gat);
not NOT_623(n2342gat,II1550);
not NOT_624(n2284gat,n2342gat);
not NOT_625(n2201gat,n2203gat);
not NOT_626(n2354gat,n2201gat);
not NOT_627(n2560gat,n2562gat);
not NOT_628(n2356gat,n2560gat);
not NOT_629(n2205gat,n2207gat);
not NOT_630(n2214gat,n2205gat);
not NOT_631(n2286gat,II1585);
not NOT_632(n2624gat,n2626gat);
not NOT_633(II1606,n2490gat);
not NOT_634(n2489gat,II1606);
not NOT_635(II1617,n2622gat);
not NOT_636(n2621gat,II1617);
not NOT_637(n2533gat,n2534gat);
not NOT_638(II1630,n2630gat);
not NOT_639(n2629gat,II1630);
not NOT_640(n2486gat,n2629gat);
not NOT_641(n2541gat,n2543gat);
not NOT_642(n2429gat,n2541gat);
not NOT_643(n2432gat,n2430gat);
not NOT_644(II1655,n2102gat);
not NOT_645(n2101gat,II1655);
not NOT_646(n1693gat,n2101gat);
not NOT_647(II1667,n1880gat);
not NOT_648(n1879gat,II1667);
not NOT_649(n1698gat,n1934gat);
not NOT_650(n1543gat,n1606gat);
not NOT_651(II1683,n1763gat);
not NOT_652(n1762gat,II1683);
not NOT_653(n1673gat,n2989gat);
not NOT_654(n1858gat,n1673gat);
not NOT_655(II1698,n2155gat);
not NOT_656(n2154gat,II1698);
not NOT_657(n2488gat,n2490gat);
not NOT_658(II1703,n2626gat);
not NOT_659(n2625gat,II1703);
not NOT_660(n2530gat,n2531gat);
not NOT_661(II1708,n2543gat);
not NOT_662(n2542gat,II1708);
not NOT_663(n2482gat,n2542gat);
not NOT_664(n2426gat,n2480gat);
not NOT_665(n2153gat,n2155gat);
not NOT_666(n2341gat,n2343gat);
not NOT_667(n2355gat,n2341gat);
not NOT_668(II1719,n2562gat);
not NOT_669(n2561gat,II1719);
not NOT_670(n2443gat,n2561gat);
not NOT_671(n2289gat,II1724);
not NOT_672(n2148gat,II1734);
not NOT_673(n855gat,n2148gat);
not NOT_674(n759gat,n855gat);
not NOT_675(II1749,n1035gat);
not NOT_676(n1034gat,II1749);
not NOT_677(II1752,n1034gat);
not NOT_678(n1189gat,II1752);
not NOT_679(n1075gat,n855gat);
not NOT_680(II1766,n1121gat);
not NOT_681(n1120gat,II1766);
not NOT_682(II1769,n1120gat);
not NOT_683(n1190gat,II1769);
not NOT_684(n760gat,n855gat);
not NOT_685(II1783,n1072gat);
not NOT_686(n1071gat,II1783);
not NOT_687(II1786,n1071gat);
not NOT_688(n1191gat,II1786);
not NOT_689(n1119gat,n1121gat);
not NOT_690(II1791,n1119gat);
not NOT_691(n1192gat,II1791);
not NOT_692(n1070gat,n1072gat);
not NOT_693(II1795,n1070gat);
not NOT_694(n1193gat,II1795);
not NOT_695(n1033gat,n1035gat);
not NOT_696(II1800,n1033gat);
not NOT_697(n1194gat,II1800);
not NOT_698(n1183gat,n1184gat);
not NOT_699(II1807,n1183gat);
not NOT_700(n1274gat,II1807);
not NOT_701(n644gat,n855gat);
not NOT_702(n1280gat,n1282gat);
not NOT_703(n641gat,n855gat);
not NOT_704(II1833,n1226gat);
not NOT_705(n1225gat,II1833);
not NOT_706(II1837,n1282gat);
not NOT_707(n1281gat,II1837);
not NOT_708(n1224gat,n1226gat);
not NOT_709(II1843,n2970gat);
not NOT_710(n1275gat,II1843);
not NOT_711(n761gat,n855gat);
not NOT_712(II1857,n931gat);
not NOT_713(n930gat,II1857);
not NOT_714(II1860,n930gat);
not NOT_715(n1206gat,II1860);
not NOT_716(n762gat,n855gat);
not NOT_717(II1874,n1135gat);
not NOT_718(n1134gat,II1874);
not NOT_719(II1877,n1134gat);
not NOT_720(n1207gat,II1877);
not NOT_721(n643gat,n855gat);
not NOT_722(II1891,n1045gat);
not NOT_723(n1044gat,II1891);
not NOT_724(II1894,n1044gat);
not NOT_725(n1208gat,II1894);
not NOT_726(n1133gat,n1135gat);
not NOT_727(II1899,n1133gat);
not NOT_728(n1209gat,II1899);
not NOT_729(n1043gat,n1045gat);
not NOT_730(II1903,n1043gat);
not NOT_731(n1210gat,II1903);
not NOT_732(n929gat,n931gat);
not NOT_733(II1908,n929gat);
not NOT_734(n1211gat,II1908);
not NOT_735(n1268gat,n1201gat);
not NOT_736(II1915,n1268gat);
not NOT_737(n1276gat,II1915);
not NOT_738(n1329gat,n2970gat);
not NOT_739(II1920,n1329gat);
not NOT_740(n1277gat,II1920);
not NOT_741(II1923,n1201gat);
not NOT_742(n1278gat,II1923);
not NOT_743(II1927,n1184gat);
not NOT_744(n1279gat,II1927);
not NOT_745(n1284gat,n1269gat);
not NOT_746(n642gat,n855gat);
not NOT_747(n1195gat,n1197gat);
not NOT_748(II1947,n1197gat);
not NOT_749(n1196gat,II1947);
not NOT_750(n2516gat,n2518gat);
not NOT_751(II1961,n2516gat);
not NOT_752(n3017gat,II1961);
not NOT_753(n851gat,n853gat);
not NOT_754(n1725gat,n2148gat);
not NOT_755(n664gat,n1725gat);
not NOT_756(n852gat,n854gat);
not NOT_757(II1981,n667gat);
not NOT_758(n666gat,II1981);
not NOT_759(n368gat,n1725gat);
not NOT_760(II1996,n659gat);
not NOT_761(n658gat,II1996);
not NOT_762(II1999,n658gat);
not NOT_763(n784gat,II1999);
not NOT_764(n662gat,n1725gat);
not NOT_765(II2014,n553gat);
not NOT_766(n552gat,II2014);
not NOT_767(II2017,n552gat);
not NOT_768(n785gat,II2017);
not NOT_769(n661gat,n1725gat);
not NOT_770(II2032,n777gat);
not NOT_771(n776gat,II2032);
not NOT_772(II2035,n776gat);
not NOT_773(n786gat,II2035);
not NOT_774(n551gat,n553gat);
not NOT_775(II2040,n551gat);
not NOT_776(n787gat,II2040);
not NOT_777(n775gat,n777gat);
not NOT_778(II2044,n775gat);
not NOT_779(n788gat,II2044);
not NOT_780(n657gat,n659gat);
not NOT_781(II2049,n657gat);
not NOT_782(n789gat,II2049);
not NOT_783(n35gat,n779gat);
not NOT_784(II2056,n35gat);
not NOT_785(n125gat,II2056);
not NOT_786(n558gat,n1725gat);
not NOT_787(n559gat,n561gat);
not NOT_788(n371gat,n1725gat);
not NOT_789(II2084,n366gat);
not NOT_790(n365gat,II2084);
not NOT_791(II2088,n561gat);
not NOT_792(n560gat,II2088);
not NOT_793(n364gat,n366gat);
not NOT_794(II2094,n2876gat);
not NOT_795(n126gat,II2094);
not NOT_796(n663gat,n1725gat);
not NOT_797(II2109,n322gat);
not NOT_798(n321gat,II2109);
not NOT_799(II2112,n321gat);
not NOT_800(n226gat,II2112);
not NOT_801(n370gat,n1725gat);
not NOT_802(II2127,n318gat);
not NOT_803(n317gat,II2127);
not NOT_804(II2130,n317gat);
not NOT_805(n227gat,II2130);
not NOT_806(n369gat,n1725gat);
not NOT_807(II2145,n314gat);
not NOT_808(n313gat,II2145);
not NOT_809(II2148,n313gat);
not NOT_810(n228gat,II2148);
not NOT_811(n316gat,n318gat);
not NOT_812(II2153,n316gat);
not NOT_813(n229gat,II2153);
not NOT_814(n312gat,n314gat);
not NOT_815(II2157,n312gat);
not NOT_816(n230gat,II2157);
not NOT_817(n320gat,n322gat);
not NOT_818(II2162,n320gat);
not NOT_819(n231gat,II2162);
not NOT_820(n34gat,n221gat);
not NOT_821(II2169,n34gat);
not NOT_822(n127gat,II2169);
not NOT_823(n133gat,n2876gat);
not NOT_824(II2174,n133gat);
not NOT_825(n128gat,II2174);
not NOT_826(II2177,n221gat);
not NOT_827(n129gat,II2177);
not NOT_828(II2181,n779gat);
not NOT_829(n130gat,II2181);
not NOT_830(n665gat,n667gat);
not NOT_831(n1601gat,n120gat);
not NOT_832(n2597gat,n2599gat);
not NOT_833(n2595gat,n2594gat);
not NOT_834(n2586gat,n2588gat);
not NOT_835(II2213,n2342gat);
not NOT_836(n2573gat,II2213);
not NOT_837(n2638gat,n2640gat);
not NOT_838(II2225,n2638gat);
not NOT_839(n2574gat,II2225);
not NOT_840(II2228,n2561gat);
not NOT_841(n2575gat,II2228);
not NOT_842(II2232,n2640gat);
not NOT_843(n2639gat,II2232);
not NOT_844(II2235,n2639gat);
not NOT_845(n2576gat,II2235);
not NOT_846(II2238,n2560gat);
not NOT_847(n2577gat,II2238);
not NOT_848(II2242,n2341gat);
not NOT_849(n2578gat,II2242);
not NOT_850(II2248,n2568gat);
not NOT_851(n2582gat,II2248);
not NOT_852(II2251,n2207gat);
not NOT_853(n2206gat,II2251);
not NOT_854(II2254,n2206gat);
not NOT_855(n2414gat,II2254);
not NOT_856(II2257,n2398gat);
not NOT_857(n2415gat,II2257);
not NOT_858(II2260,n2203gat);
not NOT_859(n2202gat,II2260);
not NOT_860(II2263,n2202gat);
not NOT_861(n2416gat,II2263);
not NOT_862(n2397gat,n2399gat);
not NOT_863(II2268,n2397gat);
not NOT_864(n2417gat,II2268);
not NOT_865(II2271,n2201gat);
not NOT_866(n2418gat,II2271);
not NOT_867(II2275,n2205gat);
not NOT_868(n2419gat,II2275);
not NOT_869(II2281,n2409gat);
not NOT_870(n2585gat,II2281);
not NOT_871(n2656gat,n2658gat);
not NOT_872(n2493gat,n2495gat);
not NOT_873(n2388gat,n2390gat);
not NOT_874(II2316,n2390gat);
not NOT_875(n2389gat,II2316);
not NOT_876(II2319,n2495gat);
not NOT_877(n2494gat,II2319);
not NOT_878(II2324,n3014gat);
not NOT_879(n2649gat,II2324);
not NOT_880(n2268gat,n2270gat);
not NOT_881(II2344,n2339gat);
not NOT_882(n2338gat,II2344);
not NOT_883(n2337gat,n2339gat);
not NOT_884(II2349,n2270gat);
not NOT_885(n2269gat,II2349);
not NOT_886(II2354,n2880gat);
not NOT_887(n2652gat,II2354);
not NOT_888(n2500gat,n2502gat);
not NOT_889(n2620gat,n2622gat);
not NOT_890(n2612gat,n2620gat);
not NOT_891(II2372,n2612gat);
not NOT_892(n2606gat,II2372);
not NOT_893(n2532gat,n2625gat);
not NOT_894(II2376,n2532gat);
not NOT_895(n2607gat,II2376);
not NOT_896(n2540gat,n2488gat);
not NOT_897(II2380,n2540gat);
not NOT_898(n2608gat,II2380);
not NOT_899(n2536gat,n2624gat);
not NOT_900(II2385,n2536gat);
not NOT_901(n2609gat,II2385);
not NOT_902(n2487gat,n2489gat);
not NOT_903(II2389,n2487gat);
not NOT_904(n2610gat,II2389);
not NOT_905(n2557gat,n2621gat);
not NOT_906(II2394,n2557gat);
not NOT_907(n2611gat,II2394);
not NOT_908(II2400,n2601gat);
not NOT_909(n2616gat,II2400);
not NOT_910(II2403,n2629gat);
not NOT_911(n2550gat,II2403);
not NOT_912(II2414,n2634gat);
not NOT_913(n2633gat,II2414);
not NOT_914(II2417,n2633gat);
not NOT_915(n2551gat,II2417);
not NOT_916(II2420,n2542gat);
not NOT_917(n2552gat,II2420);
not NOT_918(n2632gat,n2634gat);
not NOT_919(II2425,n2632gat);
not NOT_920(n2553gat,II2425);
not NOT_921(II2428,n2541gat);
not NOT_922(n2554gat,II2428);
not NOT_923(n2628gat,n2630gat);
not NOT_924(II2433,n2628gat);
not NOT_925(n2555gat,II2433);
not NOT_926(II2439,n2545gat);
not NOT_927(n2619gat,II2439);
not NOT_928(n2504gat,n2506gat);
not NOT_929(n2660gat,n2655gat);
not NOT_930(n1528gat,n2293gat);
not NOT_931(n1523gat,n2219gat);
not NOT_932(n1592gat,n1529gat);
not NOT_933(n2666gat,n1704gat);
not NOT_934(n2422gat,n3013gat);
not NOT_935(n2290gat,n2202gat);
not NOT_936(n2081gat,n2218gat);
not NOT_937(n2285gat,n2397gat);
not NOT_938(n2359gat,n2358gat);
not NOT_939(n1414gat,n1415gat);
not NOT_940(n566gat,n364gat);
not NOT_941(n1480gat,n2292gat);
not NOT_942(n1301gat,n1416gat);
not NOT_943(n1150gat,n312gat);
not NOT_944(n873gat,n316gat);
not NOT_945(n2011gat,n2306gat);
not NOT_946(n1478gat,n1481gat);
not NOT_947(n875gat,n559gat);
not NOT_948(n1410gat,n2357gat);
not NOT_949(n876gat,n1347gat);
not NOT_950(n1160gat,n1484gat);
not NOT_951(n1084gat,n657gat);
not NOT_952(n983gat,n320gat);
not NOT_953(n1482gat,n2363gat);
not NOT_954(n1157gat,n1483gat);
not NOT_955(n985gat,n775gat);
not NOT_956(n1530gat,n2364gat);
not NOT_957(n1307gat,n1308gat);
not NOT_958(n1085gat,n551gat);
not NOT_959(n1479gat,n2291gat);
not NOT_960(n1348gat,n1349gat);
not NOT_961(n2217gat,n2206gat);
not NOT_962(n1591gat,n2223gat);
not NOT_963(n1437gat,n1438gat);
not NOT_964(n1832gat,n1834gat);
not NOT_965(n1765gat,n1767gat);
not NOT_966(n1878gat,n1880gat);
not NOT_967(n1442gat,n1831gat);
not NOT_968(n1444gat,n1442gat);
not NOT_969(n1378gat,n2975gat);
not NOT_970(n1322gat,n2974gat);
not NOT_971(n1439gat,n1486gat);
not NOT_972(n1370gat,n1426gat);
not NOT_973(n1369gat,n2966gat);
not NOT_974(n1366gat,n1365gat);
not NOT_975(n1374gat,n2979gat);
not NOT_976(n2162gat,n2220gat);
not NOT_977(n1450gat,n1423gat);
not NOT_978(n1427gat,n1608gat);
not NOT_979(n1603gat,n1831gat);
not NOT_980(n2082gat,n2084gat);
not NOT_981(n1449gat,n1494gat);
not NOT_982(n1590gat,n1603gat);
not NOT_983(n1248gat,n2954gat);
not NOT_984(n1418gat,n1417gat);
not NOT_985(n1306gat,n2964gat);
not NOT_986(n1353gat,n1419gat);
not NOT_987(n1247gat,n2958gat);
not NOT_988(n1355gat,n1422gat);
not NOT_989(n1300gat,n2963gat);
not NOT_990(n1487gat,n1485gat);
not NOT_991(n1164gat,n2953gat);
not NOT_992(n1356gat,n1354gat);
not NOT_993(n1436gat,n1435gat);
not NOT_994(n1106gat,n2949gat);
not NOT_995(n1425gat,n1421gat);
not NOT_996(n1105gat,n2934gat);
not NOT_997(n1424gat,n1420gat);
not NOT_998(n1309gat,n2959gat);
not NOT_999(II2672,n2143gat);
not NOT_1000(n2142gat,II2672);
not NOT_1001(n1788gat,n2142gat);
not NOT_1002(II2684,n2061gat);
not NOT_1003(n2060gat,II2684);
not NOT_1004(n1786gat,n2060gat);
not NOT_1005(II2696,n2139gat);
not NOT_1006(n2138gat,II2696);
not NOT_1007(n1839gat,n2138gat);
not NOT_1008(n1897gat,n1899gat);
not NOT_1009(n1884gat,n1897gat);
not NOT_1010(n1848gat,n1850gat);
not NOT_1011(n1783gat,n1848gat);
not NOT_1012(n1548gat,II2721);
not NOT_1013(n1719gat,n1548gat);
not NOT_1014(n2137gat,n2139gat);
not NOT_1015(n1633gat,n2137gat);
not NOT_1016(n2059gat,n2061gat);
not NOT_1017(n1785gat,n2059gat);
not NOT_1018(II2731,n1850gat);
not NOT_1019(n1849gat,II2731);
not NOT_1020(n1784gat,n1849gat);
not NOT_1021(n1716gat,II2736);
not NOT_1022(n1635gat,n1716gat);
not NOT_1023(n2401gat,n2403gat);
not NOT_1024(n1989gat,n2401gat);
not NOT_1025(n2392gat,n2394gat);
not NOT_1026(n1918gat,n2392gat);
not NOT_1027(II2771,n2440gat);
not NOT_1028(n2439gat,II2771);
not NOT_1029(n1986gat,n2439gat);
not NOT_1030(n1866gat,n1865gat);
not NOT_1031(II2785,n2407gat);
not NOT_1032(n2406gat,II2785);
not NOT_1033(n2216gat,n2406gat);
not NOT_1034(n2345gat,n2347gat);
not NOT_1035(n1988gat,n2345gat);
not NOT_1036(n1735gat,n1861gat);
not NOT_1037(n1387gat,n1389gat);
not NOT_1038(n1694gat,II2813);
not NOT_1039(n1777gat,n1694gat);
not NOT_1040(n1781gat,n1780gat);
not NOT_1041(n2019gat,n2021gat);
not NOT_1042(n1549gat,II2832);
not NOT_1043(n1551gat,n1549gat);
not NOT_1044(II2837,n2347gat);
not NOT_1045(n2346gat,II2837);
not NOT_1046(n2152gat,n2346gat);
not NOT_1047(n2405gat,n2407gat);
not NOT_1048(n2351gat,n2405gat);
not NOT_1049(II2843,n2403gat);
not NOT_1050(n2402gat,II2843);
not NOT_1051(n2212gat,n2402gat);
not NOT_1052(II2847,n2394gat);
not NOT_1053(n2393gat,II2847);
not NOT_1054(n1991gat,n2393gat);
not NOT_1055(n1665gat,n1666gat);
not NOT_1056(n1517gat,n1578gat);
not NOT_1057(n1392gat,n1394gat);
not NOT_1058(II2873,n1496gat);
not NOT_1059(n1495gat,II2873);
not NOT_1060(n1685gat,n1604gat);
not NOT_1061(II2885,n2091gat);
not NOT_1062(n2090gat,II2885);
not NOT_1063(n1550gat,II2890);
not NOT_1064(n1552gat,n1550gat);
not NOT_1065(n1330gat,n1332gat);
not NOT_1066(n1738gat,n1740gat);
not NOT_1067(II2915,n1740gat);
not NOT_1068(n1739gat,II2915);
not NOT_1069(n1925gat,n1920gat);
not NOT_1070(n1917gat,n1921gat);
not NOT_1071(n2141gat,n2143gat);
not NOT_1072(n1787gat,n2141gat);
not NOT_1073(n1717gat,II2926);
not NOT_1074(n1859gat,n1717gat);
not NOT_1075(n1922gat,n1798gat);
not NOT_1076(n1713gat,II2935);
not NOT_1077(n1743gat,n1713gat);
not NOT_1078(n1923gat,n1864gat);
not NOT_1079(n1945gat,n1690gat);
not NOT_1080(II2953,n2179gat);
not NOT_1081(n2178gat,II2953);
not NOT_1082(n1661gat,n1660gat);
not NOT_1083(n1572gat,n1576gat);
not NOT_1084(n2438gat,n2440gat);
not NOT_1085(n2283gat,n2438gat);
not NOT_1086(n1520gat,n1582gat);
not NOT_1087(n1580gat,n1577gat);
not NOT_1088(n1990gat,n2988gat);
not NOT_1089(II2978,n2190gat);
not NOT_1090(n2189gat,II2978);
not NOT_1091(II2989,n2135gat);
not NOT_1092(n2134gat,II2989);
not NOT_1093(II3000,n2262gat);
not NOT_1094(n2261gat,II3000);
not NOT_1095(n2128gat,n2129gat);
not NOT_1096(n1836gat,n1695gat);
not NOT_1097(II3016,n2182gat);
not NOT_1098(n2181gat,II3016);
not NOT_1099(n1431gat,n1433gat);
not NOT_1100(n1314gat,n1316gat);
not NOT_1101(n1361gat,n1363gat);
not NOT_1102(II3056,n1312gat);
not NOT_1103(n1311gat,II3056);
not NOT_1104(n1707gat,n1626gat);
not NOT_1105(n1773gat,n1775gat);
not NOT_1106(n1659gat,n2987gat);
not NOT_1107(n1515gat,n1521gat);
not NOT_1108(n1736gat,n1737gat);
not NOT_1109(n1658gat,n2216gat);
not NOT_1110(n1724gat,n1732gat);
not NOT_1111(n1662gat,n1663gat);
not NOT_1112(n1656gat,n1655gat);
not NOT_1113(n1670gat,n1667gat);
not NOT_1114(n1569gat,n1570gat);
not NOT_1115(n1568gat,n1575gat);
not NOT_1116(n1727gat,n1728gat);
not NOT_1117(n1797gat,n1801gat);
not NOT_1118(n1730gat,n1731gat);
not NOT_1119(n1561gat,n1571gat);
not NOT_1120(n1668gat,n1734gat);
not NOT_1121(n1742gat,n2216gat);
not NOT_1122(n1671gat,n1669gat);
not NOT_1123(n1652gat,n1657gat);
not NOT_1124(n1648gat,n1729gat);
not NOT_1125(n1790gat,n1726gat);
not NOT_1126(n2004gat,n1929gat);
not NOT_1127(n1869gat,n1871gat);
not NOT_1128(II3143,n2592gat);
not NOT_1129(n2591gat,II3143);
not NOT_1130(n1584gat,n2989gat);
not NOT_1131(n1714gat,II3149);
not NOT_1132(n1718gat,n1714gat);
not NOT_1133(II3163,n1508gat);
not NOT_1134(n1507gat,II3163);
not NOT_1135(n1396gat,n1401gat);
not NOT_1136(II3168,n1394gat);
not NOT_1137(n1393gat,II3168);
not NOT_1138(n1409gat,n1476gat);
not NOT_1139(II3174,n1899gat);
not NOT_1140(n1898gat,II3174);
not NOT_1141(n1838gat,n1898gat);
not NOT_1142(n1712gat,II3179);
not NOT_1143(II3191,n1678gat);
not NOT_1144(n1677gat,II3191);
not NOT_1145(n2000gat,n1412gat);
not NOT_1146(n2001gat,n1412gat);
not NOT_1147(n1999gat,n2001gat);
not NOT_1148(n2307gat,n2309gat);
not NOT_1149(II3211,n2663gat);
not NOT_1150(n3018gat,II3211);
not NOT_1151(n2448gat,n2450gat);
not NOT_1152(n2661gat,n2662gat);
not NOT_1153(n2444gat,n2446gat);
not NOT_1154(II3235,n2238gat);
not NOT_1155(n3019gat,II3235);
not NOT_1156(n1310gat,n1312gat);
not NOT_1157(n199gat,n87gat);
not NOT_1158(n195gat,n184gat);
not NOT_1159(n827gat,n204gat);
not NOT_1160(n2093gat,n2095gat);
not NOT_1161(n2174gat,n2176gat);
not NOT_1162(II3273,n2169gat);
not NOT_1163(n2168gat,II3273);
not NOT_1164(n2452gat,n2454gat);
not NOT_1165(n1691gat,n2452gat);
not NOT_1166(II3287,n1691gat);
not NOT_1167(n3020gat,II3287);
not NOT_1168(II3290,n1691gat);
not NOT_1169(n3021gat,II3290);
not NOT_1170(II3293,n1691gat);
not NOT_1171(n3022gat,II3293);
not NOT_1172(n1699gat,n2452gat);
not NOT_1173(II3297,n1699gat);
not NOT_1174(n3023gat,II3297);
not NOT_1175(II3300,n1699gat);
not NOT_1176(n3024gat,II3300);
not NOT_1177(II3303,n1691gat);
not NOT_1178(n3025gat,II3303);
not NOT_1179(II3306,n1699gat);
not NOT_1180(n3026gat,II3306);
not NOT_1181(II3309,n1699gat);
not NOT_1182(n3027gat,II3309);
not NOT_1183(II3312,n1699gat);
not NOT_1184(n3028gat,II3312);
not NOT_1185(II3315,n1869gat);
not NOT_1186(n3029gat,II3315);
not NOT_1187(II3318,n1869gat);
not NOT_1188(n3030gat,II3318);
not NOT_1189(n2260gat,n2262gat);
not NOT_1190(n2257gat,n2189gat);
not NOT_1191(n2188gat,n2190gat);
not NOT_1192(n2187gat,n3004gat);
not NOT_1193(II3336,n2040gat);
not NOT_1194(n2039gat,II3336);
not NOT_1195(II3339,n1775gat);
not NOT_1196(n1774gat,II3339);
not NOT_1197(II3342,n1316gat);
not NOT_1198(n1315gat,II3342);
not NOT_1199(n2042gat,n2044gat);
not NOT_1200(n2035gat,n2037gat);
not NOT_1201(n2023gat,n2025gat);
not NOT_1202(n2097gat,n2099gat);
not NOT_1203(n1855gat,n2014gat);
not NOT_1204(II3387,n2194gat);
not NOT_1205(n3031gat,II3387);
not NOT_1206(II3390,n2261gat);
not NOT_1207(n3032gat,II3390);
not NOT_1208(n2256gat,n3032gat);
not NOT_1209(II3394,n2260gat);
not NOT_1210(n3033gat,II3394);
not NOT_1211(n2251gat,n3033gat);
not NOT_1212(n2184gat,n3003gat);
not NOT_1213(II3401,n2192gat);
not NOT_1214(n3034gat,II3401);
not NOT_1215(n2133gat,n2135gat);
not NOT_1216(n2131gat,n2185gat);
not NOT_1217(n2049gat,n3001gat);
not NOT_1218(II3412,n2057gat);
not NOT_1219(n3035gat,II3412);
not NOT_1220(n2253gat,n2189gat);
not NOT_1221(n2252gat,n2260gat);
not NOT_1222(n2248gat,n3006gat);
not NOT_1223(n2264gat,n2266gat);
not NOT_1224(II3429,n2266gat);
not NOT_1225(n2265gat,II3429);
not NOT_1226(n2492gat,n2329gat);
not NOT_1227(II3436,n2492gat);
not NOT_1228(n3036gat,II3436);
not NOT_1229(n1709gat,n1849gat);
not NOT_1230(n1845gat,n2141gat);
not NOT_1231(n1891gat,n2059gat);
not NOT_1232(n1963gat,n2137gat);
not NOT_1233(n1886gat,n1897gat);
not NOT_1234(n1968gat,n1958gat);
not NOT_1235(n1629gat,n1895gat);
not NOT_1236(n1631gat,n1848gat);
not NOT_1237(n1711gat,n2990gat);
not NOT_1238(n2200gat,n2078gat);
not NOT_1239(n2437gat,n2195gat);
not NOT_1240(II3457,n2556gat);
not NOT_1241(n3037gat,II3457);
not NOT_1242(n1956gat,n1898gat);
not NOT_1243(II3461,n1956gat);
not NOT_1244(n3038gat,II3461);
not NOT_1245(n1954gat,n3038gat);
not NOT_1246(II3465,n1886gat);
not NOT_1247(n3039gat,II3465);
not NOT_1248(n1888gat,n3039gat);
not NOT_1249(n2048gat,n2994gat);
not NOT_1250(II3472,n2539gat);
not NOT_1251(n3040gat,II3472);
not NOT_1252(n1969gat,n2142gat);
not NOT_1253(n1893gat,n2060gat);
not NOT_1254(n1892gat,n2993gat);
not NOT_1255(II3483,n2436gat);
not NOT_1256(n3041gat,II3483);
not NOT_1257(n2056gat,n2998gat);
not NOT_1258(II3491,n2387gat);
not NOT_1259(n3042gat,II3491);
not NOT_1260(II3494,n1963gat);
not NOT_1261(n3043gat,II3494);
not NOT_1262(n1960gat,n3043gat);
not NOT_1263(n1887gat,n2138gat);
not NOT_1264(n1961gat,n2996gat);
not NOT_1265(II3504,n2330gat);
not NOT_1266(n3044gat,II3504);
not NOT_1267(n2199gat,n2147gat);
not NOT_1268(II3509,n2438gat);
not NOT_1269(n3045gat,II3509);
not NOT_1270(n2332gat,n3045gat);
not NOT_1271(II3513,n2439gat);
not NOT_1272(n3046gat,II3513);
not NOT_1273(n2259gat,n3046gat);
not NOT_1274(n2328gat,n3008gat);
not NOT_1275(II3520,n2498gat);
not NOT_1276(n3047gat,II3520);
not NOT_1277(n2151gat,n2193gat);
not NOT_1278(n2209gat,n3005gat);
not NOT_1279(II3530,n2396gat);
not NOT_1280(n3048gat,II3530);
not NOT_1281(n2052gat,n2393gat);
not NOT_1282(n2058gat,n2997gat);
not NOT_1283(II3539,n2198gat);
not NOT_1284(n3049gat,II3539);
not NOT_1285(n2349gat,n2215gat);
not NOT_1286(n2281gat,n3009gat);
not NOT_1287(II3549,n2197gat);
not NOT_1288(n3050gat,II3549);
not NOT_1289(n2146gat,n3002gat);
not NOT_1290(II3558,n2196gat);
not NOT_1291(n3051gat,II3558);
not NOT_1292(n2031gat,n2033gat);
not NOT_1293(n2108gat,n2110gat);
not NOT_1294(II3587,n2125gat);
not NOT_1295(n2124gat,II3587);
not NOT_1296(n2123gat,n2125gat);
not NOT_1297(n2119gat,n2121gat);
not NOT_1298(n2115gat,n2117gat);
not NOT_1299(II3610,n1882gat);
not NOT_1300(n3052gat,II3610);
not NOT_1301(II3621,n1975gat);
not NOT_1302(n1974gat,II3621);
not NOT_1303(n1955gat,n1956gat);
not NOT_1304(n1970gat,n1896gat);
not NOT_1305(n1973gat,n1975gat);
not NOT_1306(n2558gat,n2559gat);
not NOT_1307(II3635,n2558gat);
not NOT_1308(n3053gat,II3635);
not NOT_1309(II3646,n2644gat);
not NOT_1310(n2643gat,II3646);
not NOT_1311(n2333gat,n2438gat);
not NOT_1312(n2564gat,n2352gat);
not NOT_1313(n2642gat,n2644gat);
not NOT_1314(n2636gat,n2637gat);
not NOT_1315(II3660,n2636gat);
not NOT_1316(n3054gat,II3660);
not NOT_1317(n88gat,n84gat);
not NOT_1318(n375gat,n110gat);
not NOT_1319(II3677,n156gat);
not NOT_1320(n155gat,II3677);
not NOT_1321(n253gat,n1702gat);
not NOT_1322(n150gat,n152gat);
not NOT_1323(II3691,n152gat);
not NOT_1324(n151gat,II3691);
not NOT_1325(n243gat,n1702gat);
not NOT_1326(n233gat,n243gat);
not NOT_1327(n154gat,n156gat);
not NOT_1328(n800gat,n2874gat);
not NOT_1329(II3703,n2917gat);
not NOT_1330(n3055gat,II3703);
not NOT_1331(n235gat,n2878gat);
not NOT_1332(II3713,n2892gat);
not NOT_1333(n3056gat,II3713);
not NOT_1334(n372gat,n212gat);
not NOT_1335(n329gat,n331gat);
not NOT_1336(II3736,n388gat);
not NOT_1337(n387gat,II3736);
not NOT_1338(n334gat,n1700gat);
not NOT_1339(n386gat,n388gat);
not NOT_1340(II3742,n331gat);
not NOT_1341(n330gat,II3742);
not NOT_1342(n1430gat,n1700gat);
not NOT_1343(n1490gat,n1430gat);
not NOT_1344(n452gat,n2885gat);
not NOT_1345(II3754,n2900gat);
not NOT_1346(n3057gat,II3754);
not NOT_1347(n333gat,n2883gat);
not NOT_1348(II3765,n2929gat);
not NOT_1349(n3058gat,II3765);
not NOT_1350(II3777,n463gat);
not NOT_1351(n462gat,II3777);
not NOT_1352(n325gat,n327gat);
not NOT_1353(n457gat,n2884gat);
not NOT_1354(n461gat,n463gat);
not NOT_1355(n458gat,n2902gat);
not NOT_1356(II3801,n2925gat);
not NOT_1357(n3059gat,II3801);
not NOT_1358(n144gat,n247gat);
not NOT_1359(II3808,n327gat);
not NOT_1360(n326gat,II3808);
not NOT_1361(n878gat,n2879gat);
not NOT_1362(II3817,n2916gat);
not NOT_1363(n3060gat,II3817);
not NOT_1364(n382gat,n384gat);
not NOT_1365(II3831,n384gat);
not NOT_1366(n383gat,II3831);
not NOT_1367(n134gat,n2875gat);
not NOT_1368(II3841,n2899gat);
not NOT_1369(n3061gat,II3841);
not NOT_1370(n254gat,n256gat);
not NOT_1371(n252gat,n2877gat);
not NOT_1372(n468gat,n470gat);
not NOT_1373(II3867,n470gat);
not NOT_1374(n469gat,II3867);
not NOT_1375(n381gat,n2893gat);
not NOT_1376(II3876,n2926gat);
not NOT_1377(n3062gat,II3876);
not NOT_1378(n241gat,n140gat);
not NOT_1379(II3882,n256gat);
not NOT_1380(n255gat,II3882);
not NOT_1381(n802gat,n2882gat);
not NOT_1382(II3891,n2924gat);
not NOT_1383(n3063gat,II3891);
not NOT_1384(n146gat,n148gat);
not NOT_1385(II3904,n148gat);
not NOT_1386(n147gat,II3904);
not NOT_1387(n380gat,n2881gat);
not NOT_1388(II3914,n2923gat);
not NOT_1389(n3064gat,II3914);
not NOT_1390(n69gat,n68gat);
not NOT_1391(n1885gat,n2048gat);
not NOT_1392(II3923,n2710gat);
not NOT_1393(n2707gat,II3923);
not NOT_1394(n16gat,n564gat);
not NOT_1395(n295gat,n357gat);
not NOT_1396(n11gat,n12gat);
not NOT_1397(n1889gat,n1961gat);
not NOT_1398(II3935,n2704gat);
not NOT_1399(n2700gat,II3935);
not NOT_1400(n2051gat,n2056gat);
not NOT_1401(II3941,n2684gat);
not NOT_1402(n2680gat,II3941);
not NOT_1403(n1350gat,n1831gat);
not NOT_1404(II3945,n1350gat);
not NOT_1405(n2696gat,II3945);
not NOT_1406(II3948,n2696gat);
not NOT_1407(n2692gat,II3948);
not NOT_1408(II3951,n2448gat);
not NOT_1409(n2683gat,II3951);
not NOT_1410(II3954,n2683gat);
not NOT_1411(n2679gat,II3954);
not NOT_1412(II3957,n2450gat);
not NOT_1413(n2449gat,II3957);
not NOT_1414(n1754gat,n2449gat);
not NOT_1415(II3962,n2830gat);
not NOT_1416(n2827gat,II3962);
not NOT_1417(n2590gat,n2592gat);
not NOT_1418(n2456gat,n2458gat);
not NOT_1419(n2512gat,n2514gat);
not NOT_1420(n1544gat,n1625gat);
not NOT_1421(n1769gat,n1771gat);
not NOT_1422(n1683gat,n1756gat);
not NOT_1423(n2167gat,n2169gat);
not NOT_1424(n2013gat,II4000);
not NOT_1425(n1791gat,n2013gat);
not NOT_1426(n2691gat,n2695gat);
not NOT_1427(n1518gat,n1694gat);
not NOT_1428(n2699gat,n2703gat);
not NOT_1429(n2159gat,n1412gat);
not NOT_1430(n2478gat,n2579gat);
not NOT_1431(II4014,n2744gat);
not NOT_1432(n2740gat,II4014);
not NOT_1433(n2158gat,n1412gat);
not NOT_1434(n2186gat,n2613gat);
not NOT_1435(II4020,n2800gat);
not NOT_1436(n2797gat,II4020);
not NOT_1437(n2288gat,II4024);
not NOT_1438(n1513gat,n2288gat);
not NOT_1439(n2537gat,n2538gat);
not NOT_1440(n2442gat,n2483gat);
not NOT_1441(n1334gat,n1336gat);
not NOT_1442(II4055,n1748gat);
not NOT_1443(n1747gat,II4055);
not NOT_1444(II4067,n1675gat);
not NOT_1445(n1674gat,II4067);
not NOT_1446(n1403gat,n1402gat);
not NOT_1447(II4081,n1807gat);
not NOT_1448(n1806gat,II4081);
not NOT_1449(n1634gat,n1712gat);
not NOT_1450(n1338gat,n1340gat);
not NOT_1451(II4105,n1456gat);
not NOT_1452(n1455gat,II4105);
not NOT_1453(II4108,n1340gat);
not NOT_1454(n1339gat,II4108);
not NOT_1455(n1505gat,n2980gat);
not NOT_1456(II4117,n1505gat);
not NOT_1457(n2758gat,II4117);
not NOT_1458(n2755gat,n2758gat);
not NOT_1459(n1546gat,n2980gat);
not NOT_1460(II4122,n1546gat);
not NOT_1461(n2752gat,II4122);
not NOT_1462(n2748gat,n2752gat);
not NOT_1463(n2012gat,n2016gat);
not NOT_1464(n2002gat,n2008gat);
not NOT_1465(II4129,n3097gat);
not NOT_1466(n2858gat,II4129);
not NOT_1467(n2857gat,n2858gat);
not NOT_1468(II4135,n3098gat);
not NOT_1469(n2766gat,II4135);
not NOT_1470(II4138,n2766gat);
not NOT_1471(n2765gat,II4138);
not NOT_1472(n1684gat,n1759gat);
not NOT_1473(n1632gat,II4145);
not NOT_1474(II4157,n1525gat);
not NOT_1475(n1524gat,II4157);
not NOT_1476(n1862gat,n1863gat);
not NOT_1477(n1919gat,n1860gat);
not NOT_1478(n1460gat,n1462gat);
not NOT_1479(II4185,n1596gat);
not NOT_1480(n1595gat,II4185);
not NOT_1481(n1454gat,n1469gat);
not NOT_1482(n1468gat,n1519gat);
not NOT_1483(II4194,n1462gat);
not NOT_1484(n1461gat,II4194);
not NOT_1485(n1477gat,n2984gat);
not NOT_1486(n1594gat,n1596gat);
not NOT_1487(II4212,n1588gat);
not NOT_1488(n1587gat,II4212);
not NOT_1489(n1681gat,II4217);
not NOT_1490(II4222,n1761gat);
not NOT_1491(n2751gat,II4222);
not NOT_1492(n2747gat,n2751gat);
not NOT_1493(II4227,n1760gat);
not NOT_1494(n2743gat,II4227);
not NOT_1495(n2739gat,n2743gat);
not NOT_1496(n1978gat,n2286gat);
not NOT_1497(II4233,n1721gat);
not NOT_1498(n2808gat,II4233);
not NOT_1499(II4236,n2808gat);
not NOT_1500(n2804gat,II4236);
not NOT_1501(n517gat,n518gat);
not NOT_1502(n417gat,n418gat);
not NOT_1503(n413gat,n411gat);
not NOT_1504(n412gat,n522gat);
not NOT_1505(n406gat,n516gat);
not NOT_1506(n407gat,n355gat);
not NOT_1507(n290gat,n525gat);
not NOT_1508(n527gat,n356gat);
not NOT_1509(n416gat,n415gat);
not NOT_1510(n528gat,n521gat);
not NOT_1511(n358gat,n532gat);
not NOT_1512(n639gat,n523gat);
not NOT_1513(n1111gat,n635gat);
not NOT_1514(n524gat,n414gat);
not NOT_1515(n1112gat,n630gat);
not NOT_1516(n741gat,n629gat);
not NOT_1517(n633gat,n634gat);
not NOT_1518(n926gat,n632gat);
not NOT_1519(n670gat,n636gat);
not NOT_1520(n1123gat,n632gat);
not NOT_1521(n1007gat,n635gat);
not NOT_1522(n1006gat,n630gat);
not NOT_1523(II4309,n2941gat);
not NOT_1524(n2814gat,II4309);
not NOT_1525(II4312,n2814gat);
not NOT_1526(n2811gat,II4312);
not NOT_1527(n1002gat,n2946gat);
not NOT_1528(II4329,n2950gat);
not NOT_1529(n2813gat,II4329);
not NOT_1530(II4332,n2813gat);
not NOT_1531(n2810gat,II4332);
not NOT_1532(n888gat,n2933gat);
not NOT_1533(II4349,n2935gat);
not NOT_1534(n2818gat,II4349);
not NOT_1535(II4352,n2818gat);
not NOT_1536(n2816gat,II4352);
not NOT_1537(n898gat,n2940gat);
not NOT_1538(II4369,n2937gat);
not NOT_1539(n2817gat,II4369);
not NOT_1540(II4372,n2817gat);
not NOT_1541(n2815gat,II4372);
not NOT_1542(n1179gat,n2947gat);
not NOT_1543(II4389,n2956gat);
not NOT_1544(n2824gat,II4389);
not NOT_1545(II4392,n2824gat);
not NOT_1546(n2821gat,II4392);
not NOT_1547(n897gat,n2939gat);
not NOT_1548(II4409,n2938gat);
not NOT_1549(n2823gat,II4409);
not NOT_1550(II4412,n2823gat);
not NOT_1551(n2820gat,II4412);
not NOT_1552(n894gat,n2932gat);
not NOT_1553(II4429,n2936gat);
not NOT_1554(n2829gat,II4429);
not NOT_1555(II4432,n2829gat);
not NOT_1556(n2826gat,II4432);
not NOT_1557(n1180gat,n2948gat);
not NOT_1558(II4449,n2955gat);
not NOT_1559(n2828gat,II4449);
not NOT_1560(II4452,n2828gat);
not NOT_1561(n2825gat,II4452);
not NOT_1562(n671gat,n673gat);
not NOT_1563(n628gat,n631gat);
not NOT_1564(n976gat,n628gat);
not NOT_1565(II4475,n2951gat);
not NOT_1566(n2807gat,II4475);
not NOT_1567(II4478,n2807gat);
not NOT_1568(n2803gat,II4478);
not NOT_1569(n2127gat,n2389gat);
not NOT_1570(II4482,n2127gat);
not NOT_1571(n2682gat,II4482);
not NOT_1572(II4485,n2682gat);
not NOT_1573(n2678gat,II4485);
not NOT_1574(n2046gat,n2269gat);
not NOT_1575(II4489,n2046gat);
not NOT_1576(n2681gat,II4489);
not NOT_1577(II4492,n2681gat);
not NOT_1578(n2677gat,II4492);
not NOT_1579(n1708gat,n2338gat);
not NOT_1580(II4496,n1708gat);
not NOT_1581(n2688gat,II4496);
not NOT_1582(II4499,n2688gat);
not NOT_1583(n2686gat,II4499);
not NOT_1584(n455gat,n291gat);
not NOT_1585(n2237gat,n2646gat);
not NOT_1586(II4506,n2764gat);
not NOT_1587(n2763gat,II4506);
not NOT_1588(n1782gat,n2971gat);
not NOT_1589(II4512,n2762gat);
not NOT_1590(n2760gat,II4512);
not NOT_1591(n2325gat,n3010gat);
not NOT_1592(II4518,n2761gat);
not NOT_1593(n2759gat,II4518);
not NOT_1594(n2245gat,n504gat);
not NOT_1595(II4524,n2757gat);
not NOT_1596(n2754gat,II4524);
not NOT_1597(n2244gat,n567gat);
not NOT_1598(II4530,n2756gat);
not NOT_1599(n2753gat,II4530);
not NOT_1600(n2243gat,n55gat);
not NOT_1601(II4536,n2750gat);
not NOT_1602(n2746gat,II4536);
not NOT_1603(n2246gat,n933gat);
not NOT_1604(II4542,n2749gat);
not NOT_1605(n2745gat,II4542);
not NOT_1606(n2384gat,n43gat);
not NOT_1607(II4548,n2742gat);
not NOT_1608(n2738gat,II4548);
not NOT_1609(n2385gat,n748gat);
not NOT_1610(II4554,n2741gat);
not NOT_1611(n2737gat,II4554);
not NOT_1612(n1286gat,n1269gat);
not NOT_1613(II4558,n1286gat);
not NOT_1614(n2687gat,II4558);
not NOT_1615(n2685gat,n2687gat);
not NOT_1616(n1328gat,n1224gat);
not NOT_1617(n1381gat,n1328gat);
not NOT_1618(n1384gat,n2184gat);
not NOT_1619(II4566,n2694gat);
not NOT_1620(n2690gat,II4566);
not NOT_1621(n1382gat,n1280gat);
not NOT_1622(n1451gat,n1382gat);
not NOT_1623(n1453gat,n2187gat);
not NOT_1624(II4573,n2693gat);
not NOT_1625(n2689gat,II4573);
not NOT_1626(n927gat,n1133gat);
not NOT_1627(n925gat,n927gat);
not NOT_1628(n1452gat,n2049gat);
not NOT_1629(II4580,n2702gat);
not NOT_1630(n2698gat,II4580);
not NOT_1631(n923gat,n1043gat);
not NOT_1632(n921gat,n923gat);
not NOT_1633(n1890gat,n2328gat);
not NOT_1634(II4587,n2701gat);
not NOT_1635(n2697gat,II4587);
not NOT_1636(n850gat,n929gat);
not NOT_1637(n739gat,n850gat);
not NOT_1638(n1841gat,n2058gat);
not NOT_1639(II4594,n2709gat);
not NOT_1640(n2706gat,II4594);
not NOT_1641(n922gat,n1119gat);
not NOT_1642(n848gat,n922gat);
not NOT_1643(n2047gat,n2209gat);
not NOT_1644(II4601,n2708gat);
not NOT_1645(n2705gat,II4601);
not NOT_1646(n924gat,n1070gat);
not NOT_1647(n849gat,n924gat);
not NOT_1648(n2050gat,n2146gat);
not NOT_1649(II4608,n2799gat);
not NOT_1650(n2796gat,II4608);
not NOT_1651(n1118gat,n1033gat);
not NOT_1652(n1032gat,n1118gat);
not NOT_1653(n2054gat,n2281gat);
not NOT_1654(II4615,n2798gat);
not NOT_1655(n2795gat,II4615);
not NOT_1656(II4620,n1745gat);
not NOT_1657(n2806gat,II4620);
not NOT_1658(II4623,n2806gat);
not NOT_1659(n2802gat,II4623);
not NOT_1660(II4626,n1871gat);
not NOT_1661(n1870gat,II4626);
not NOT_1662(n1086gat,n1870gat);
not NOT_1663(II4630,n1086gat);
not NOT_1664(n2805gat,II4630);
not NOT_1665(II4633,n2805gat);
not NOT_1666(n2801gat,II4633);
not NOT_1667(n67gat,n85gat);
not NOT_1668(n71gat,n180gat);
not NOT_1669(n1840gat,n1892gat);
not NOT_1670(II4642,n2812gat);
not NOT_1671(n2809gat,II4642);
not NOT_1672(n76gat,n82gat);
not NOT_1673(n14gat,n186gat);
not NOT_1674(n1842gat,n1711gat);
not NOT_1675(II4651,n2822gat);
not NOT_1676(n2819gat,II4651);
not NOT_1677(II4654,n2819gat);
not NOT_1678(n3104gat,II4654);
not NOT_1679(II4657,n2809gat);
not NOT_1680(n3105gat,II4657);
not NOT_1681(II4660,n2801gat);
not NOT_1682(n3106gat,II4660);
not NOT_1683(II4663,n2802gat);
not NOT_1684(n3107gat,II4663);
not NOT_1685(II4666,n2795gat);
not NOT_1686(n3108gat,II4666);
not NOT_1687(II4669,n2796gat);
not NOT_1688(n3109gat,II4669);
not NOT_1689(II4672,n2705gat);
not NOT_1690(n3110gat,II4672);
not NOT_1691(II4675,n2706gat);
not NOT_1692(n3111gat,II4675);
not NOT_1693(II4678,n2697gat);
not NOT_1694(n3112gat,II4678);
not NOT_1695(II4681,n2698gat);
not NOT_1696(n3113gat,II4681);
not NOT_1697(II4684,n2689gat);
not NOT_1698(n3114gat,II4684);
not NOT_1699(II4687,n2690gat);
not NOT_1700(n3115gat,II4687);
not NOT_1701(II4690,n2685gat);
not NOT_1702(n3116gat,II4690);
not NOT_1703(II4693,n2737gat);
not NOT_1704(n3117gat,II4693);
not NOT_1705(II4696,n2738gat);
not NOT_1706(n3118gat,II4696);
not NOT_1707(II4699,n2745gat);
not NOT_1708(n3119gat,II4699);
not NOT_1709(II4702,n2746gat);
not NOT_1710(n3120gat,II4702);
not NOT_1711(II4705,n2753gat);
not NOT_1712(n3121gat,II4705);
not NOT_1713(II4708,n2754gat);
not NOT_1714(n3122gat,II4708);
not NOT_1715(II4711,n2759gat);
not NOT_1716(n3123gat,II4711);
not NOT_1717(II4714,n2760gat);
not NOT_1718(n3124gat,II4714);
not NOT_1719(II4717,n2763gat);
not NOT_1720(n3125gat,II4717);
not NOT_1721(II4720,n2686gat);
not NOT_1722(n3126gat,II4720);
not NOT_1723(II4723,n2677gat);
not NOT_1724(n3127gat,II4723);
not NOT_1725(II4726,n2678gat);
not NOT_1726(n3128gat,II4726);
not NOT_1727(II4729,n2803gat);
not NOT_1728(n3129gat,II4729);
not NOT_1729(II4732,n2825gat);
not NOT_1730(n3130gat,II4732);
not NOT_1731(II4735,n2826gat);
not NOT_1732(n3131gat,II4735);
not NOT_1733(II4738,n2820gat);
not NOT_1734(n3132gat,II4738);
not NOT_1735(II4741,n2821gat);
not NOT_1736(n3133gat,II4741);
not NOT_1737(II4744,n2815gat);
not NOT_1738(n3134gat,II4744);
not NOT_1739(II4747,n2816gat);
not NOT_1740(n3135gat,II4747);
not NOT_1741(II4750,n2810gat);
not NOT_1742(n3136gat,II4750);
not NOT_1743(II4753,n2811gat);
not NOT_1744(n3137gat,II4753);
not NOT_1745(II4756,n2804gat);
not NOT_1746(n3138gat,II4756);
not NOT_1747(II4759,n2739gat);
not NOT_1748(n3139gat,II4759);
not NOT_1749(II4762,n2747gat);
not NOT_1750(n3140gat,II4762);
not NOT_1751(II4765,n2748gat);
not NOT_1752(n3141gat,II4765);
not NOT_1753(II4768,n2755gat);
not NOT_1754(n3142gat,II4768);
not NOT_1755(II4771,n2797gat);
not NOT_1756(n3143gat,II4771);
not NOT_1757(II4774,n2740gat);
not NOT_1758(n3144gat,II4774);
not NOT_1759(II4777,n2699gat);
not NOT_1760(n3145gat,II4777);
not NOT_1761(II4780,n2691gat);
not NOT_1762(n3146gat,II4780);
not NOT_1763(II4783,n2827gat);
not NOT_1764(n3147gat,II4783);
not NOT_1765(II4786,n2679gat);
not NOT_1766(n3148gat,II4786);
not NOT_1767(II4789,n2692gat);
not NOT_1768(n3149gat,II4789);
not NOT_1769(II4792,n2680gat);
not NOT_1770(n3150gat,II4792);
not NOT_1771(II4795,n2700gat);
not NOT_1772(n3151gat,II4795);
not NOT_1773(II4798,n2707gat);
not NOT_1774(n3152gat,II4798);
or OR2_0(n2897gat,n648gat,n442gat);
or OR4_0(n1213gat,n1214gat,n1215gat,n1216gat,n1217gat);
or OR2_1(n2906gat,n745gat,n638gat);
or OR2_2(n2889gat,n423gat,n362gat);
or OR4_1(n748gat,n749gat,n750gat,n751gat,n752gat);
or OR4_2(n258gat,n259gat,n260gat,n261gat,n262gat);
or OR4_3(n1013gat,n1014gat,n1015gat,n1016gat,n1017gat);
or OR4_4(n475gat,n476gat,n477gat,n478gat,n479gat);
or OR4_5(n43gat,n44gat,n45gat,n46gat,n47gat);
or OR2_3(n2786gat,n3091gat,n3092gat);
or OR4_6(n167gat,n168gat,n169gat,n170gat,n171gat);
or OR4_7(n906gat,n907gat,n908gat,n909gat,n910gat);
or OR4_8(n343gat,n344gat,n345gat,n346gat,n347gat);
or OR4_9(n55gat,n56gat,n57gat,n58gat,n59gat);
or OR2_4(n2914gat,n768gat,n655gat);
or OR2_5(n2928gat,n963gat,n868gat);
or OR2_6(n2927gat,n962gat,n959gat);
or OR4_10(n944gat,n945gat,n946gat,n947gat,n948gat);
or OR2_7(n2896gat,n647gat,n441gat);
or OR2_8(n2922gat,n967gat,n792gat);
or OR4_11(n1228gat,n1229gat,n1230gat,n1231gat,n1232gat);
or OR2_9(n2894gat,n443gat,n439gat);
or OR2_10(n2921gat,n966gat,n790gat);
or OR2_11(n2895gat,n444gat,n440gat);
or OR4_12(n1050gat,n1051gat,n1052gat,n1053gat,n1054gat);
or OR4_13(n933gat,n934gat,n935gat,n936gat,n937gat);
or OR4_14(n709gat,n710gat,n711gat,n712gat,n713gat);
or OR4_15(n728gat,n729gat,n730gat,n731gat,n732gat);
or OR4_16(n493gat,n494gat,n495gat,n496gat,n497gat);
or OR4_17(n504gat,n505gat,n506gat,n507gat,n508gat);
or OR3_0(II1277,n2860gat,n2855gat,n2863gat);
or OR3_1(II1278,n740gat,n3030gat,II1277);
or OR2_12(n2913gat,n767gat,n653gat);
or OR2_13(n2920gat,n867gat,n771gat);
or OR2_14(n2905gat,n964gat,n961gat);
or OR4_18(n803gat,n804gat,n805gat,n806gat,n807gat);
or OR4_19(n586gat,n587gat,n588gat,n589gat,n590gat);
or OR2_15(n2898gat,n447gat,n445gat);
or OR4_20(n686gat,n687gat,n688gat,n689gat,n690gat);
or OR4_21(n567gat,n568gat,n569gat,n570gat,n571gat);
or OR3_2(II1515,n2474gat,n2524gat,n2831gat);
or OR3_3(II1516,n2466gat,n2462gat,II1515);
or OR3_4(II1584,n2353gat,n2284gat,n2354gat);
or OR3_5(II1585,n2356gat,n2214gat,II1584);
or OR2_16(n2989gat,n1693gat,n1692gat);
or OR3_6(II1723,n2354gat,n2353gat,n2214gat);
or OR3_7(II1724,n2355gat,n2443gat,II1723);
or OR3_8(II1733,n2286gat,n2428gat,n2289gat);
or OR3_9(II1734,n1604gat,n2214gat,II1733);
or OR2_17(n2918gat,n769gat,n759gat);
or OR2_18(n2952gat,n1076gat,n1075gat);
or OR2_19(n2919gat,n766gat,n760gat);
or OR4_22(n1184gat,n1185gat,n1186gat,n1187gat,n1188gat);
or OR2_20(n2910gat,n645gat,n644gat);
or OR2_21(n2907gat,n646gat,n641gat);
or OR2_22(n2970gat,n1383gat,n1327gat);
or OR2_23(n2911gat,n761gat,n651gat);
or OR2_24(n2912gat,n762gat,n652gat);
or OR2_25(n2909gat,n765gat,n643gat);
or OR4_23(n1201gat,n1202gat,n1203gat,n1204gat,n1205gat);
or OR4_24(n1269gat,n1270gat,n1271gat,n1272gat,n1273gat);
or OR2_26(n2908gat,n763gat,n642gat);
or OR2_27(n2971gat,n1287gat,n1285gat);
or OR3_10(n2904gat,n793gat,n664gat,n556gat);
or OR3_11(n2891gat,n795gat,n656gat,n368gat);
or OR3_12(n2903gat,n794gat,n773gat,n662gat);
or OR3_13(n2915gat,n965gat,n960gat,n661gat);
or OR4_25(n779gat,n780gat,n781gat,n782gat,n783gat);
or OR3_14(n2901gat,n558gat,n555gat,n450gat);
or OR3_15(n2890gat,n654gat,n557gat,n371gat);
or OR2_28(n2876gat,n874gat,n132gat);
or OR3_16(n2888gat,n663gat,n649gat,n449gat);
or OR3_17(n2887gat,n791gat,n650gat,n370gat);
or OR3_18(n2886gat,n774gat,n764gat,n369gat);
or OR4_26(n221gat,n222gat,n223gat,n224gat,n225gat);
or OR4_27(n120gat,n121gat,n122gat,n123gat,n124gat);
or OR2_29(n3010gat,n2460gat,n2423gat);
or OR2_30(n3016gat,n2596gat,n2595gat);
or OR4_28(n2568gat,n2569gat,n2570gat,n2571gat,n2572gat);
or OR4_29(n2409gat,n2410gat,n2411gat,n2412gat,n2413gat);
or OR2_31(n2579gat,n2580gat,n2581gat);
or OR2_32(n3014gat,n2567gat,n2499gat);
or OR2_33(n2880gat,n299gat,n207gat);
or OR2_34(n2646gat,n2647gat,n2648gat);
or OR4_30(n2601gat,n2602gat,n2603gat,n2604gat,n2605gat);
or OR4_31(n2545gat,n2546gat,n2547gat,n2548gat,n2549gat);
or OR2_35(n2613gat,n2614gat,n2615gat);
or OR2_36(n3013gat,n2461gat,n2421gat);
or OR4_32(n2930gat,n1153gat,n1151gat,n982gat,n877gat);
or OR4_33(n2957gat,n1159gat,n1158gat,n1156gat,n1155gat);
or OR2_37(n2975gat,n1443gat,n1325gat);
or OR2_38(n2974gat,n1321gat,n1320gat);
or OR2_39(n2966gat,n1368gat,n1258gat);
or OR2_40(n2979gat,n1373gat,n1372gat);
or OR4_34(n2978gat,n1441gat,n1440gat,n1371gat,n1367gat);
or OR2_41(n2982gat,n1504gat,n1502gat);
or OR2_42(n2954gat,n1250gat,n1103gat);
or OR2_43(n2964gat,n1304gat,n1249gat);
or OR2_44(n2958gat,n1246gat,n1161gat);
or OR2_45(n2963gat,n1291gat,n1245gat);
or OR4_35(n2973gat,n1352gat,n1351gat,n1303gat,n1302gat);
or OR2_46(n2953gat,n1163gat,n1102gat);
or OR2_47(n2949gat,n1101gat,n996gat);
or OR2_48(n2934gat,n1104gat,n887gat);
or OR2_49(n2959gat,n1305gat,n1162gat);
or OR4_36(n2977gat,n1360gat,n1359gat,n1358gat,n1357gat);
or OR3_19(II2720,n1788gat,n1786gat,n1839gat);
or OR3_20(II2721,n1884gat,n1783gat,II2720);
or OR3_21(II2735,n1788gat,n1884gat,n1633gat);
or OR3_22(II2736,n1785gat,n1784gat,II2735);
or OR3_23(II2812,n1703gat,n1704gat,n1778gat);
or OR4_37(II2813,n1609gat,n1702gat,n1700gat,II2812);
or OR3_24(II2831,n1839gat,n1786gat,n1788gat);
or OR3_25(II2832,n1884gat,n1784gat,II2831);
or OR3_26(II2889,n1784gat,n1633gat,n1884gat);
or OR3_27(II2890,n1788gat,n1786gat,II2889);
or OR3_28(II2925,n1784gat,n1785gat,n1633gat);
or OR3_29(II2926,n1884gat,n1787gat,II2925);
or OR3_30(II2934,n1784gat,n1839gat,n1788gat);
or OR3_31(II2935,n1785gat,n1884gat,II2934);
or OR2_50(n2988gat,n1733gat,n1581gat);
or OR2_51(n2983gat,n2079gat,n2073gat);
or OR2_52(n2987gat,n1574gat,n1573gat);
or OR3_32(n2992gat,n1723gat,n1647gat,n1646gat);
or OR3_33(n2986gat,n1650gat,n1649gat,n1563gat);
or OR3_34(n2991gat,n1654gat,n1653gat,n1644gat);
or OR3_35(II3148,n1839gat,n1884gat,n1784gat);
or OR3_36(II3149,n1786gat,n1787gat,II3148);
or OR3_37(II3178,n1838gat,n1785gat,n1788gat);
or OR3_38(II3179,n1839gat,n1784gat,II3178);
or OR3_39(n2981gat,n1413gat,n1408gat,n1407gat);
or OR2_53(n3000gat,n2000gat,n1999gat);
or OR3_40(n3004gat,n2258gat,n2257gat,n2255gat);
or OR2_54(n3003gat,n2256gat,n2251gat);
or OR2_55(n3001gat,n2132gat,n2130gat);
or OR2_56(n3006gat,n2253gat,n2252gat);
or OR2_57(n3007gat,n2250gat,n2249gat);
or OR2_58(n2990gat,n1710gat,n1630gat);
or OR2_59(n2994gat,n1954gat,n1888gat);
or OR3_41(n2993gat,n1894gat,n1847gat,n1846gat);
or OR2_60(n2998gat,n2055gat,n1967gat);
or OR3_42(n2996gat,n1960gat,n1959gat,n1957gat);
or OR2_61(n3008gat,n2332gat,n2259gat);
or OR2_62(n3005gat,n2211gat,n2210gat);
or OR3_43(n2997gat,n2053gat,n2052gat,n1964gat);
or OR2_63(n3009gat,n2350gat,n2282gat);
or OR3_44(n3002gat,n2213gat,n2150gat,n2149gat);
or OR2_64(n2995gat,n1962gat,n1955gat);
or OR2_65(n2999gat,n1972gat,n1971gat);
or OR2_66(n3011gat,n2333gat,n2331gat);
or OR2_67(n3015gat,n2566gat,n2565gat);
or OR3_45(n2874gat,n141gat,n38gat,n37gat);
or OR2_68(n2917gat,n1074gat,n872gat);
or OR2_69(n2878gat,n234gat,n137gat);
or OR2_70(n2892gat,n378gat,n377gat);
or OR3_46(n2885gat,n250gat,n249gat,n248gat);
or OR3_47(n2900gat,n869gat,n453gat,n448gat);
or OR2_71(n2883gat,n251gat,n244gat);
or OR3_48(n2929gat,n974gat,n973gat,n870gat);
or OR2_72(n2884gat,n246gat,n245gat);
or OR2_73(n2902gat,n460gat,n459gat);
or OR3_49(n2925gat,n975gat,n972gat,n969gat);
or OR2_74(n2879gat,n145gat,n143gat);
or OR3_50(n2916gat,n971gat,n970gat,n968gat);
or OR3_51(n2875gat,n142gat,n40gat,n39gat);
or OR3_52(n2899gat,n772gat,n451gat,n446gat);
or OR2_75(n2877gat,n139gat,n136gat);
or OR2_76(n2893gat,n391gat,n390gat);
or OR2_77(n2926gat,n1083gat,n1077gat);
or OR2_78(n2882gat,n242gat,n240gat);
or OR2_79(n2924gat,n871gat,n797gat);
or OR3_53(n2881gat,n324gat,n238gat,n237gat);
or OR2_80(n2923gat,n1082gat,n796gat);
or OR2_81(n2710gat,n69gat,n1885gat);
or OR2_82(n2704gat,n11gat,n1889gat);
or OR2_83(n2684gat,n1599gat,n2051gat);
or OR2_84(n2830gat,n2444gat,n1754gat);
or OR3_54(II3999,n2167gat,n2031gat,n2174gat);
or OR4_38(II4000,n2108gat,n2093gat,n2035gat,II3999);
or OR2_85(n2695gat,n1586gat,n1791gat);
or OR2_86(n2703gat,n1755gat,n1518gat);
or OR2_87(n2744gat,n2159gat,n2478gat);
or OR2_88(n2800gat,n2158gat,n2186gat);
or OR3_55(II4023,n2443gat,n2290gat,n2214gat);
or OR3_56(II4024,n2353gat,n2284gat,II4023);
or OR4_39(n2980gat,n1470gat,n1400gat,n1399gat,n1398gat);
or OR3_57(II4144,n1633gat,n1838gat,n1786gat);
or OR3_58(II4145,n1788gat,n1784gat,II4144);
or OR2_89(n2984gat,n1467gat,n1466gat);
or OR4_40(n2985gat,n1686gat,n1533gat,n1532gat,n1531gat);
or OR3_59(II4216,n1427gat,n1595gat,n1677gat);
or OR3_60(II4217,n1392gat,n2989gat,II4216);
or OR4_41(n2931gat,n1100gat,n994gat,n989gat,n880gat);
or OR2_90(n2943gat,n1012gat,n905gat);
or OR2_91(n2941gat,n1003gat,n902gat);
or OR4_42(n2946gat,n1099gat,n998gat,n995gat,n980gat);
or OR2_92(n2960gat,n1175gat,n1174gat);
or OR2_93(n2950gat,n1001gat,n999gat);
or OR2_94(n2969gat,n1323gat,n1264gat);
or OR4_43(n2933gat,n981gat,n890gat,n889gat,n886gat);
or OR2_95(n2935gat,n892gat,n891gat);
or OR2_96(n2942gat,n904gat,n903gat);
or OR4_44(n2940gat,n1152gat,n1092gat,n997gat,n993gat);
or OR2_97(n2937gat,n900gat,n895gat);
or OR4_45(n2947gat,n1094gat,n1093gat,n988gat,n984gat);
or OR2_98(n2965gat,n1267gat,n1257gat);
or OR2_99(n2956gat,n1178gat,n1116gat);
or OR2_100(n2961gat,n1375gat,n1324gat);
or OR4_46(n2939gat,n1091gat,n1088gat,n992gat,n987gat);
or OR2_101(n2938gat,n899gat,n896gat);
or OR2_102(n2967gat,n1262gat,n1260gat);
or OR4_47(n2932gat,n1098gat,n1090gat,n986gat,n885gat);
or OR2_103(n2936gat,n901gat,n893gat);
or OR4_48(n2948gat,n1097gat,n1089gat,n1087gat,n991gat);
or OR2_104(n2968gat,n1326gat,n1261gat);
or OR2_105(n2955gat,n1177gat,n1115gat);
or OR2_106(n2944gat,n977gat,n976gat);
or OR4_49(n2945gat,n1096gat,n1095gat,n990gat,n979gat);
or OR2_107(n2962gat,n1176gat,n1173gat);
or OR2_108(n2951gat,n1004gat,n1000gat);
or OR2_109(n2764gat,n1029gat,n2237gat);
or OR2_110(n2762gat,n1028gat,n1782gat);
or OR2_111(n2761gat,n1031gat,n2325gat);
or OR2_112(n2757gat,n1030gat,n2245gat);
or OR2_113(n2756gat,n1011gat,n2244gat);
or OR2_114(n2750gat,n1181gat,n2243gat);
or OR2_115(n2749gat,n1010gat,n2246gat);
or OR2_116(n2742gat,n1005gat,n2384gat);
or OR2_117(n2741gat,n1182gat,n2385gat);
or OR2_118(n2694gat,n1381gat,n1384gat);
or OR2_119(n2693gat,n1451gat,n1453gat);
or OR2_120(n2702gat,n925gat,n1452gat);
or OR2_121(n2701gat,n921gat,n1890gat);
or OR2_122(n2709gat,n739gat,n1841gat);
or OR2_123(n2708gat,n848gat,n2047gat);
or OR2_124(n2799gat,n849gat,n2050gat);
or OR2_125(n2798gat,n1032gat,n2054gat);
or OR3_61(n2812gat,n73gat,n70gat,n1840gat);
or OR3_62(n2822gat,n77gat,n13gat,n1842gat);
nor NOR2_0(n421gat,n2715gat,n2723gat);
nor NOR2_1(n648gat,n373gat,n2669gat);
nor NOR2_2(n442gat,n2844gat,n856gat);
nor NOR2_3(n1499gat,n396gat,n401gat);
nor NOR2_4(n1616gat,n918gat,n396gat);
nor NOR2_5(n1614gat,n396gat,n845gat);
nor NOR3_0(n1641gat,n1645gat,n1553gat,n1559gat);
nor NOR3_1(n1642gat,n1559gat,n1616gat,n1645gat);
nor NOR3_2(n1556gat,n1614gat,n1645gat,n1616gat);
nor NOR3_3(n1557gat,n1553gat,n1645gat,n1614gat);
nor NOR3_4(n1639gat,n1499gat,n1559gat,n1553gat);
nor NOR4_0(n1605gat,n1614gat,n1616gat,n1499gat,n396gat);
nor NOR3_5(n1555gat,n1616gat,n1559gat,n1499gat);
nor NOR3_6(n1558gat,n1614gat,n1553gat,n1499gat);
nor NOR2_6(n1256gat,n392gat,n702gat);
nor NOR2_7(n1117gat,n720gat,n725gat);
nor NOR2_8(n1618gat,n1319gat,n1447gat);
nor NOR2_9(n1114gat,n725gat,n721gat);
nor NOR2_10(n1621gat,n1319gat,n1380gat);
nor NOR2_11(n1318gat,n392gat,n701gat);
nor NOR2_12(n1619gat,n1447gat,n1446gat);
nor NOR2_13(n1622gat,n1380gat,n1446gat);
nor NOR3_7(n1214gat,n1218gat,n1219gat,n1220gat);
nor NOR3_8(n1215gat,n1218gat,n1221gat,n1222gat);
nor NOR3_9(n1216gat,n1223gat,n1219gat,n1222gat);
nor NOR3_10(n1217gat,n1223gat,n1221gat,n1220gat);
nor NOR2_14(n745gat,n2716gat,n2867gat);
nor NOR2_15(n638gat,n2715gat,n2868gat);
nor NOR2_16(n423gat,n2724gat,n2726gat);
nor NOR2_17(n362gat,n2723gat,n2727gat);
nor NOR3_11(n749gat,n753gat,n754gat,n755gat);
nor NOR3_12(n750gat,n753gat,n756gat,n757gat);
nor NOR3_13(n751gat,n758gat,n754gat,n757gat);
nor NOR3_14(n752gat,n758gat,n756gat,n755gat);
nor NOR3_15(n259gat,n263gat,n264gat,n265gat);
nor NOR3_16(n260gat,n263gat,n266gat,n267gat);
nor NOR3_17(n261gat,n268gat,n264gat,n267gat);
nor NOR3_18(n262gat,n268gat,n266gat,n265gat);
nor NOR3_19(n1014gat,n1018gat,n1019gat,n1020gat);
nor NOR3_20(n1015gat,n1018gat,n1021gat,n1022gat);
nor NOR3_21(n1016gat,n1023gat,n1019gat,n1022gat);
nor NOR3_22(n1017gat,n1023gat,n1021gat,n1020gat);
nor NOR3_23(n476gat,n480gat,n481gat,n482gat);
nor NOR3_24(n477gat,n480gat,n483gat,n484gat);
nor NOR3_25(n478gat,n485gat,n481gat,n484gat);
nor NOR3_26(n479gat,n485gat,n483gat,n482gat);
nor NOR3_27(n44gat,n48gat,n49gat,n50gat);
nor NOR3_28(n45gat,n48gat,n51gat,n52gat);
nor NOR3_29(n46gat,n53gat,n49gat,n52gat);
nor NOR3_30(n47gat,n53gat,n51gat,n50gat);
nor NOR2_18(n1376gat,n724gat,n720gat);
nor NOR2_19(n1617gat,n1319gat,n1448gat);
nor NOR2_20(n1377gat,n724gat,n721gat);
nor NOR2_21(n1624gat,n1319gat,n1379gat);
nor NOR2_22(n1113gat,n393gat,n701gat);
nor NOR2_23(n1501gat,n1448gat,n1500gat);
nor NOR2_24(n1623gat,n1379gat,n1446gat);
nor NOR2_25(n1620gat,n1448gat,n1446gat);
nor NOR2_26(n1827gat,n2729gat,n2317gat);
nor NOR2_27(n1817gat,n1819gat,n1823gat);
nor NOR2_28(n1935gat,n1816gat,n1828gat);
nor NOR2_29(n529gat,n2724gat,n2715gat);
nor NOR2_30(n361gat,n2859gat,n2726gat);
nor NOR3_31(n168gat,n172gat,n173gat,n174gat);
nor NOR3_32(n169gat,n172gat,n175gat,n176gat);
nor NOR3_33(n170gat,n177gat,n173gat,n176gat);
nor NOR3_34(n171gat,n177gat,n175gat,n174gat);
nor NOR3_35(n907gat,n911gat,n912gat,n913gat);
nor NOR3_36(n908gat,n911gat,n914gat,n915gat);
nor NOR3_37(n909gat,n916gat,n912gat,n915gat);
nor NOR3_38(n910gat,n916gat,n914gat,n913gat);
nor NOR3_39(n344gat,n348gat,n349gat,n350gat);
nor NOR3_40(n345gat,n348gat,n351gat,n352gat);
nor NOR3_41(n346gat,n353gat,n349gat,n352gat);
nor NOR3_42(n347gat,n353gat,n351gat,n350gat);
nor NOR3_43(n56gat,n60gat,n61gat,n62gat);
nor NOR3_44(n57gat,n60gat,n63gat,n64gat);
nor NOR3_45(n58gat,n65gat,n61gat,n64gat);
nor NOR3_46(n59gat,n65gat,n63gat,n62gat);
nor NOR2_31(n768gat,n373gat,n2731gat);
nor NOR2_32(n655gat,n856gat,n2718gat);
nor NOR2_33(n963gat,n856gat,n2838gat);
nor NOR2_34(n868gat,n2775gat,n373gat);
nor NOR2_35(n962gat,n856gat,n2711gat);
nor NOR2_36(n959gat,n373gat,n2734gat);
nor NOR3_47(n945gat,n949gat,n950gat,n951gat);
nor NOR3_48(n946gat,n949gat,n952gat,n953gat);
nor NOR3_49(n947gat,n954gat,n950gat,n953gat);
nor NOR3_50(n948gat,n954gat,n952gat,n951gat);
nor NOR2_37(n647gat,n2792gat,n373gat);
nor NOR2_38(n441gat,n856gat,n2846gat);
nor NOR2_39(n967gat,n373gat,n2672gat);
nor NOR2_40(n792gat,n2852gat,n856gat);
nor NOR3_51(n1229gat,n1233gat,n1234gat,n1235gat);
nor NOR3_52(n1230gat,n1233gat,n1236gat,n1237gat);
nor NOR3_53(n1231gat,n1238gat,n1234gat,n1237gat);
nor NOR3_54(n1232gat,n1238gat,n1236gat,n1235gat);
nor NOR2_41(n443gat,n2778gat,n373gat);
nor NOR2_42(n439gat,n856gat,n2836gat);
nor NOR2_43(n966gat,n2789gat,n373gat);
nor NOR2_44(n790gat,n856gat,n2840gat);
nor NOR2_45(n444gat,n373gat,n2781gat);
nor NOR2_46(n440gat,n856gat,n2842gat);
nor NOR3_55(n1051gat,n1055gat,n1056gat,n1057gat);
nor NOR3_56(n1052gat,n1055gat,n1058gat,n1059gat);
nor NOR3_57(n1053gat,n1060gat,n1056gat,n1059gat);
nor NOR3_58(n1054gat,n1060gat,n1058gat,n1057gat);
nor NOR3_59(n934gat,n938gat,n939gat,n940gat);
nor NOR3_60(n935gat,n938gat,n941gat,n942gat);
nor NOR3_61(n936gat,n943gat,n939gat,n942gat);
nor NOR3_62(n937gat,n943gat,n941gat,n940gat);
nor NOR2_47(n746gat,n2716gat,n2723gat);
nor NOR2_48(n360gat,n2859gat,n2727gat);
nor NOR3_63(n710gat,n714gat,n715gat,n716gat);
nor NOR3_64(n711gat,n714gat,n717gat,n718gat);
nor NOR3_65(n712gat,n719gat,n715gat,n718gat);
nor NOR3_66(n713gat,n719gat,n717gat,n716gat);
nor NOR3_67(n729gat,n733gat,n734gat,n735gat);
nor NOR3_68(n730gat,n733gat,n736gat,n737gat);
nor NOR3_69(n731gat,n738gat,n734gat,n737gat);
nor NOR3_70(n732gat,n738gat,n736gat,n735gat);
nor NOR3_71(n494gat,n498gat,n499gat,n500gat);
nor NOR3_72(n495gat,n498gat,n501gat,n502gat);
nor NOR3_73(n496gat,n503gat,n499gat,n502gat);
nor NOR3_74(n497gat,n503gat,n501gat,n500gat);
nor NOR3_75(n505gat,n509gat,n510gat,n511gat);
nor NOR3_76(n506gat,n509gat,n512gat,n513gat);
nor NOR3_77(n507gat,n514gat,n510gat,n513gat);
nor NOR3_78(n508gat,n514gat,n512gat,n511gat);
nor NOR4_1(n564gat,n3029gat,n2863gat,n2855gat,n374gat);
nor NOR3_79(n86gat,n743gat,n294gat,n17gat);
nor NOR2_49(n78gat,n2784gat,n79gat);
nor NOR2_50(n767gat,n219gat,n2731gat);
nor NOR2_51(n286gat,n289gat,n2723gat);
nor NOR2_52(n287gat,n289gat,n2715gat);
nor NOR2_53(n288gat,n289gat,n2726gat);
nor NOR3_80(n181gat,n286gat,n179gat,n188gat);
nor NOR2_54(n182gat,n72gat,n2720gat);
nor NOR2_55(n653gat,n2718gat,n111gat);
nor NOR2_56(n867gat,n219gat,n2775gat);
nor NOR2_57(n771gat,n2838gat,n111gat);
nor NOR2_58(n964gat,n111gat,n2711gat);
nor NOR2_59(n961gat,n219gat,n2734gat);
nor NOR3_81(n804gat,n808gat,n809gat,n810gat);
nor NOR3_82(n805gat,n808gat,n811gat,n812gat);
nor NOR3_83(n806gat,n813gat,n809gat,n812gat);
nor NOR3_84(n807gat,n813gat,n811gat,n810gat);
nor NOR3_85(n587gat,n591gat,n592gat,n593gat);
nor NOR3_86(n588gat,n591gat,n594gat,n595gat);
nor NOR3_87(n589gat,n596gat,n592gat,n595gat);
nor NOR3_88(n590gat,n596gat,n594gat,n593gat);
nor NOR2_60(n447gat,n2836gat,n111gat);
nor NOR2_61(n445gat,n2778gat,n219gat);
nor NOR3_89(n687gat,n691gat,n692gat,n693gat);
nor NOR3_90(n688gat,n691gat,n694gat,n695gat);
nor NOR3_91(n689gat,n696gat,n692gat,n695gat);
nor NOR3_92(n690gat,n696gat,n694gat,n693gat);
nor NOR3_93(n568gat,n572gat,n573gat,n574gat);
nor NOR3_94(n569gat,n572gat,n575gat,n576gat);
nor NOR3_95(n570gat,n577gat,n573gat,n576gat);
nor NOR3_96(n571gat,n577gat,n575gat,n574gat);
nor NOR3_97(n187gat,n189gat,n287gat,n188gat);
nor NOR2_62(n197gat,n194gat,n297gat);
nor NOR3_98(n15gat,n637gat,n17gat,n293gat);
nor NOR2_63(n22gat,n92gat,n21gat);
nor NOR2_64(n93gat,n197gat,n22gat);
nor NOR2_65(n769gat,n93gat,n2731gat);
nor NOR3_99(n2534gat,n2624gat,n2489gat,n2621gat);
nor NOR3_100(n2430gat,n2533gat,n2486gat,n2429gat);
nor NOR2_66(n1606gat,n3020gat,n270gat);
nor NOR2_67(n2239gat,n2850gat,n3019gat);
nor NOR3_101(n1934gat,n2470gat,n1935gat,n2239gat);
nor NOR2_68(n1610gat,n1698gat,n1543gat);
nor NOR2_69(n1692gat,n1879gat,n1762gat);
nor NOR2_70(n2433gat,n2432gat,n2154gat);
nor NOR3_102(n2531gat,n2488gat,n2625gat,n2621gat);
nor NOR3_103(n2480gat,n2530gat,n2482gat,n2486gat);
nor NOR2_71(n2427gat,n2426gat,n2153gat);
nor NOR2_72(n2428gat,n2433gat,n2427gat);
nor NOR2_73(n1778gat,n3026gat,n1779gat);
nor NOR2_74(n1609gat,n1503gat,n3025gat);
nor NOR2_75(n1702gat,n3024gat,n1615gat);
nor NOR2_76(n1700gat,n1701gat,n3023gat);
nor NOR4_2(n1604gat,n1778gat,n1609gat,n1702gat,n1700gat);
nor NOR2_77(n1076gat,n93gat,n2775gat);
nor NOR2_78(n766gat,n93gat,n2734gat);
nor NOR3_104(n1185gat,n1189gat,n1190gat,n1191gat);
nor NOR3_105(n1186gat,n1189gat,n1192gat,n1193gat);
nor NOR3_106(n1187gat,n1194gat,n1190gat,n1193gat);
nor NOR3_107(n1188gat,n1194gat,n1192gat,n1191gat);
nor NOR2_79(n645gat,n2792gat,n93gat);
nor NOR2_80(n646gat,n93gat,n2669gat);
nor NOR2_81(n1383gat,n1280gat,n1225gat);
nor NOR2_82(n1327gat,n1281gat,n1224gat);
nor NOR2_83(n651gat,n93gat,n2778gat);
nor NOR2_84(n652gat,n2789gat,n93gat);
nor NOR2_85(n765gat,n2781gat,n93gat);
nor NOR3_108(n1202gat,n1206gat,n1207gat,n1208gat);
nor NOR3_109(n1203gat,n1206gat,n1209gat,n1210gat);
nor NOR3_110(n1204gat,n1211gat,n1207gat,n1210gat);
nor NOR3_111(n1205gat,n1211gat,n1209gat,n1208gat);
nor NOR3_112(n1270gat,n1274gat,n1275gat,n1276gat);
nor NOR3_113(n1271gat,n1274gat,n1277gat,n1278gat);
nor NOR3_114(n1272gat,n1279gat,n1275gat,n1278gat);
nor NOR3_115(n1273gat,n1279gat,n1277gat,n1276gat);
nor NOR2_86(n763gat,n2672gat,n93gat);
nor NOR2_87(n1287gat,n1284gat,n1195gat);
nor NOR2_88(n1285gat,n1196gat,n1269gat);
nor NOR2_89(n853gat,n740gat,n2148gat);
nor NOR2_90(n793gat,n2852gat,n851gat);
nor NOR2_91(n854gat,n2148gat,n374gat);
nor NOR2_92(n556gat,n2672gat,n852gat);
nor NOR2_93(n795gat,n2731gat,n852gat);
nor NOR2_94(n656gat,n851gat,n2718gat);
nor NOR2_95(n794gat,n852gat,n2775gat);
nor NOR2_96(n773gat,n851gat,n2838gat);
nor NOR2_97(n965gat,n2711gat,n851gat);
nor NOR2_98(n960gat,n2734gat,n852gat);
nor NOR3_116(n780gat,n784gat,n785gat,n786gat);
nor NOR3_117(n781gat,n784gat,n787gat,n788gat);
nor NOR3_118(n782gat,n789gat,n785gat,n788gat);
nor NOR3_119(n783gat,n789gat,n787gat,n786gat);
nor NOR2_99(n555gat,n852gat,n2792gat);
nor NOR2_100(n450gat,n851gat,n2846gat);
nor NOR2_101(n654gat,n851gat,n2844gat);
nor NOR2_102(n557gat,n2669gat,n852gat);
nor NOR2_103(n874gat,n559gat,n365gat);
nor NOR2_104(n132gat,n560gat,n364gat);
nor NOR2_105(n649gat,n2778gat,n852gat);
nor NOR2_106(n449gat,n2836gat,n851gat);
nor NOR2_107(n791gat,n851gat,n2840gat);
nor NOR2_108(n650gat,n852gat,n2789gat);
nor NOR2_109(n774gat,n2842gat,n851gat);
nor NOR2_110(n764gat,n852gat,n2781gat);
nor NOR3_120(n222gat,n226gat,n227gat,n228gat);
nor NOR3_121(n223gat,n226gat,n229gat,n230gat);
nor NOR3_122(n224gat,n231gat,n227gat,n230gat);
nor NOR3_123(n225gat,n231gat,n229gat,n228gat);
nor NOR3_124(n121gat,n125gat,n126gat,n127gat);
nor NOR3_125(n122gat,n125gat,n128gat,n129gat);
nor NOR3_126(n123gat,n130gat,n126gat,n129gat);
nor NOR3_127(n124gat,n130gat,n128gat,n127gat);
nor NOR2_111(n2460gat,n666gat,n120gat);
nor NOR2_112(n2423gat,n665gat,n1601gat);
nor NOR3_128(n2594gat,n3017gat,n2520gat,n2597gat);
nor NOR3_129(n2569gat,n2573gat,n2574gat,n2575gat);
nor NOR3_130(n2570gat,n2573gat,n2576gat,n2577gat);
nor NOR3_131(n2571gat,n2578gat,n2574gat,n2577gat);
nor NOR3_132(n2572gat,n2578gat,n2576gat,n2575gat);
nor NOR3_133(n2410gat,n2414gat,n2415gat,n2416gat);
nor NOR3_134(n2411gat,n2414gat,n2417gat,n2418gat);
nor NOR3_135(n2412gat,n2419gat,n2415gat,n2418gat);
nor NOR3_136(n2413gat,n2419gat,n2417gat,n2416gat);
nor NOR2_113(n2583gat,n2582gat,n2585gat);
nor NOR2_114(n2580gat,n2582gat,n2583gat);
nor NOR2_115(n2581gat,n2583gat,n2585gat);
nor NOR2_116(n2567gat,n2493gat,n2388gat);
nor NOR2_117(n2499gat,n2389gat,n2494gat);
nor NOR2_118(n299gat,n2268gat,n2338gat);
nor NOR2_119(n207gat,n2337gat,n2269gat);
nor NOR2_120(n2650gat,n2649gat,n2652gat);
nor NOR2_121(n2647gat,n2649gat,n2650gat);
nor NOR2_122(n2648gat,n2650gat,n2652gat);
nor NOR3_137(n2602gat,n2606gat,n2607gat,n2608gat);
nor NOR3_138(n2603gat,n2606gat,n2609gat,n2610gat);
nor NOR3_139(n2604gat,n2611gat,n2607gat,n2610gat);
nor NOR3_140(n2605gat,n2611gat,n2609gat,n2608gat);
nor NOR3_141(n2546gat,n2550gat,n2551gat,n2552gat);
nor NOR3_142(n2547gat,n2550gat,n2553gat,n2554gat);
nor NOR3_143(n2548gat,n2555gat,n2551gat,n2554gat);
nor NOR3_144(n2549gat,n2555gat,n2553gat,n2552gat);
nor NOR2_123(n2617gat,n2616gat,n2619gat);
nor NOR2_124(n2614gat,n2616gat,n2617gat);
nor NOR2_125(n2615gat,n2617gat,n2619gat);
nor NOR4_3(n2655gat,n2508gat,n2656gat,n2500gat,n2504gat);
nor NOR3_145(n2293gat,n2353gat,n2284gat,n2443gat);
nor NOR2_126(n2219gat,n2354gat,n2214gat);
nor NOR2_127(n1529gat,n1528gat,n1523gat);
nor NOR2_128(n1704gat,n3027gat,n1706gat);
nor NOR2_129(n2461gat,n120gat,n2666gat);
nor NOR2_130(n2421gat,n1601gat,n1704gat);
nor NOR2_131(n1598gat,n1592gat,n2422gat);
nor NOR2_132(n2218gat,n2214gat,n2290gat);
nor NOR3_146(n2358gat,n2285gat,n2356gat,n2355gat);
nor NOR2_133(n1415gat,n2081gat,n2359gat);
nor NOR2_134(n1153gat,n1414gat,n566gat);
nor NOR3_147(n2292gat,n2443gat,n2284gat,n2285gat);
nor NOR2_135(n1416gat,n2081gat,n1480gat);
nor NOR2_136(n1151gat,n1301gat,n1150gat);
nor NOR3_148(n2306gat,n2356gat,n2284gat,n2285gat);
nor NOR2_137(n1481gat,n2081gat,n2011gat);
nor NOR2_138(n982gat,n873gat,n1478gat);
nor NOR3_149(n2357gat,n2285gat,n2355gat,n2443gat);
nor NOR2_139(n1347gat,n2081gat,n1410gat);
nor NOR2_140(n877gat,n875gat,n876gat);
nor NOR2_141(n1484gat,n2081gat,n1528gat);
nor NOR2_142(n1159gat,n1160gat,n1084gat);
nor NOR3_150(n2363gat,n2353gat,n2356gat,n2355gat);
nor NOR2_143(n1483gat,n2081gat,n1482gat);
nor NOR2_144(n1158gat,n983gat,n1157gat);
nor NOR3_151(n2364gat,n2353gat,n2284gat,n2356gat);
nor NOR2_145(n1308gat,n2081gat,n1530gat);
nor NOR2_146(n1156gat,n985gat,n1307gat);
nor NOR3_152(n2291gat,n2353gat,n2355gat,n2443gat);
nor NOR2_147(n1349gat,n1479gat,n2081gat);
nor NOR2_148(n1155gat,n1085gat,n1348gat);
nor NOR3_153(n1154gat,n1598gat,n2930gat,n2957gat);
nor NOR2_149(n1703gat,n1705gat,n3028gat);
nor NOR2_150(n1608gat,n1704gat,n1703gat);
nor NOR2_151(n1411gat,n1154gat,n1608gat);
nor NOR2_152(n2223gat,n2354gat,n2217gat);
nor NOR2_153(n1438gat,n1591gat,n1480gat);
nor NOR2_154(n1625gat,n3021gat,n1628gat);
nor NOR2_155(n1626gat,n1627gat,n3022gat);
nor NOR3_154(n1831gat,n1832gat,n1765gat,n1878gat);
nor NOR2_156(n1443gat,n1442gat,n706gat);
nor NOR2_157(n1325gat,n1444gat,n164gat);
nor NOR2_158(n1441gat,n1437gat,n1378gat);
nor NOR2_159(n1321gat,n1442gat,n837gat);
nor NOR2_160(n1320gat,n1444gat,n278gat);
nor NOR2_161(n1486gat,n1482gat,n1591gat);
nor NOR2_162(n1440gat,n1322gat,n1439gat);
nor NOR2_163(n1426gat,n2011gat,n1591gat);
nor NOR2_164(n1368gat,n1442gat,n613gat);
nor NOR2_165(n1258gat,n274gat,n1444gat);
nor NOR2_166(n1371gat,n1370gat,n1369gat);
nor NOR2_167(n1365gat,n1479gat,n1591gat);
nor NOR2_168(n1373gat,n833gat,n1442gat);
nor NOR2_169(n1372gat,n282gat,n1444gat);
nor NOR2_170(n1367gat,n1366gat,n1374gat);
nor NOR2_171(n2220gat,n2290gat,n2217gat);
nor NOR2_172(n1423gat,n2162gat,n1530gat);
nor NOR2_173(n1498gat,n1609gat,n1427gat);
nor NOR2_174(n1504gat,n1450gat,n1498gat);
nor NOR2_175(n1607gat,n2082gat,n1609gat);
nor NOR2_176(n1494gat,n1528gat,n2162gat);
nor NOR2_177(n1502gat,n1607gat,n1449gat);
nor NOR2_178(n1250gat,n1603gat,n815gat);
nor NOR2_179(n1103gat,n956gat,n1590gat);
nor NOR2_180(n1417gat,n2162gat,n1480gat);
nor NOR2_181(n1352gat,n1248gat,n1418gat);
nor NOR2_182(n1304gat,n1590gat,n1067gat);
nor NOR2_183(n1249gat,n679gat,n1603gat);
nor NOR2_184(n1419gat,n2162gat,n1479gat);
nor NOR2_185(n1351gat,n1306gat,n1353gat);
nor NOR2_186(n1246gat,n864gat,n1590gat);
nor NOR2_187(n1161gat,n583gat,n1603gat);
nor NOR2_188(n1422gat,n2011gat,n2162gat);
nor NOR2_189(n1303gat,n1247gat,n1355gat);
nor NOR2_190(n1291gat,n1603gat,n579gat);
nor NOR2_191(n1245gat,n1590gat,n860gat);
nor NOR2_192(n1485gat,n1482gat,n2162gat);
nor NOR2_193(n1302gat,n1300gat,n1487gat);
nor NOR2_194(n1163gat,n882gat,n1603gat);
nor NOR2_195(n1102gat,n1297gat,n1590gat);
nor NOR2_196(n1354gat,n1591gat,n1530gat);
nor NOR2_197(n1360gat,n1164gat,n1356gat);
nor NOR2_198(n1435gat,n1591gat,n1528gat);
nor NOR2_199(n1101gat,n1590gat,n1293gat);
nor NOR2_200(n996gat,n1603gat,n823gat);
nor NOR2_201(n1359gat,n1436gat,n1106gat);
nor NOR2_202(n1421gat,n2162gat,n2359gat);
nor NOR2_203(n1104gat,n1079gat,n1590gat);
nor NOR2_204(n887gat,n1603gat,n683gat);
nor NOR2_205(n1358gat,n1425gat,n1105gat);
nor NOR2_206(n1420gat,n1410gat,n2162gat);
nor NOR2_207(n1305gat,n1147gat,n1590gat);
nor NOR2_208(n1162gat,n698gat,n1603gat);
nor NOR2_209(n1357gat,n1424gat,n1309gat);
nor NOR4_4(n1428gat,n2978gat,n2982gat,n2973gat,n2977gat);
nor NOR2_210(n1794gat,n1673gat,n1719gat);
nor NOR2_211(n1796gat,n1858gat,n1635gat);
nor NOR2_212(n1792gat,n1794gat,n1796gat);
nor NOR3_155(n1865gat,n1989gat,n1918gat,n1986gat);
nor NOR3_156(n1861gat,n1866gat,n2216gat,n1988gat);
nor NOR2_213(n1793gat,n1792gat,n1735gat);
nor NOR2_214(n1406gat,n1428gat,n1387gat);
nor NOR3_157(n1780gat,n1777gat,n1625gat,n1626gat);
nor NOR2_215(n2016gat,n2019gat,n1878gat);
nor NOR2_216(n2664gat,n2850gat,n3018gat);
nor NOR3_158(n1666gat,n1986gat,n2212gat,n1991gat);
nor NOR3_159(n1578gat,n2152gat,n2351gat,n1665gat);
nor NOR2_217(n1516gat,n1551gat,n1517gat);
nor NOR3_160(n1864gat,n1858gat,n1495gat,n2090gat);
nor NOR2_218(n1565gat,n1735gat,n1552gat);
nor NOR2_219(n1921gat,n1738gat,n1673gat);
nor NOR2_220(n1798gat,n1739gat,n1673gat);
nor NOR3_161(n1920gat,n1864gat,n1921gat,n1798gat);
nor NOR2_221(n1926gat,n1925gat,n1635gat);
nor NOR2_222(n1916gat,n1917gat,n1859gat);
nor NOR2_223(n1994gat,n1719gat,n1922gat);
nor NOR2_224(n1924gat,n1743gat,n1923gat);
nor NOR4_5(n2078gat,n1926gat,n1916gat,n1994gat,n1924gat);
nor NOR2_225(n1690gat,n1700gat,n1702gat);
nor NOR3_162(n1660gat,n1918gat,n1986gat,n2212gat);
nor NOR3_163(n1576gat,n2351gat,n1988gat,n1661gat);
nor NOR2_226(n1733gat,n1673gat,n1572gat);
nor NOR3_164(n1582gat,n2283gat,n1991gat,n2212gat);
nor NOR3_165(n1577gat,n1520gat,n2351gat,n1988gat);
nor NOR2_227(n1581gat,n1858gat,n1580gat);
nor NOR3_166(n2129gat,n2189gat,n2134gat,n2261gat);
nor NOR4_6(n2079gat,n2078gat,n2178gat,n1990gat,n2128gat);
nor NOR4_7(n1695gat,n1609gat,n1778gat,n1704gat,n1703gat);
nor NOR3_167(n2073gat,n2078gat,n1990gat,n2181gat);
nor NOR2_228(n1696gat,n1707gat,n1698gat);
nor NOR2_229(n1758gat,n1311gat,n1773gat);
nor NOR3_168(n1574gat,n1719gat,n1673gat,n1444gat);
nor NOR3_169(n1573gat,n1444gat,n1858gat,n1635gat);
nor NOR2_230(n1521gat,n2283gat,n1991gat);
nor NOR2_231(n1737gat,n2212gat,n2152gat);
nor NOR3_170(n1732gat,n1515gat,n1736gat,n1658gat);
nor NOR3_171(n1723gat,n1659gat,n1722gat,n1724gat);
nor NOR2_232(n1663gat,n1986gat,n1918gat);
nor NOR3_172(n1655gat,n1736gat,n1662gat,n1658gat);
nor NOR3_173(n1647gat,n1656gat,n1659gat,n1554gat);
nor NOR2_233(n1667gat,n1991gat,n1986gat);
nor NOR3_174(n1570gat,n1736gat,n1658gat,n1670gat);
nor NOR3_175(n1646gat,n1569gat,n1659gat,n1566gat);
nor NOR2_234(n1575gat,n1918gat,n2283gat);
nor NOR3_176(n1728gat,n1568gat,n1736gat,n1658gat);
nor NOR3_177(n1650gat,n1727gat,n1659gat,n1640gat);
nor NOR2_235(n1801gat,n2152gat,n1989gat);
nor NOR3_178(n1731gat,n1658gat,n1515gat,n1797gat);
nor NOR3_179(n1649gat,n1560gat,n1659gat,n1730gat);
nor NOR3_180(n1571gat,n1670gat,n1658gat,n1797gat);
nor NOR3_181(n1563gat,n1561gat,n1562gat,n1659gat);
nor NOR2_236(n1734gat,n1988gat,n2212gat);
nor NOR3_182(n1669gat,n1668gat,n1742gat,n1670gat);
nor NOR2_237(n1654gat,n1671gat,n1659gat);
nor NOR3_183(n1657gat,n1662gat,n1797gat,n1658gat);
nor NOR3_184(n1653gat,n1651gat,n1652gat,n1659gat);
nor NOR3_185(n1729gat,n1658gat,n1797gat,n1568gat);
nor NOR3_186(n1644gat,n1643gat,n1648gat,n1659gat);
nor NOR3_187(n1726gat,n2992gat,n2986gat,n2991gat);
nor NOR2_238(n1929gat,n1758gat,n1790gat);
nor NOR3_188(n2009gat,n2016gat,n2664gat,n2004gat);
nor NOR3_189(n1413gat,n1869gat,n672gat,n2591gat);
nor NOR2_239(n1636gat,n1584gat,n1718gat);
nor NOR2_240(n1401gat,n1584gat,n1590gat);
nor NOR3_190(n1408gat,n1507gat,n1396gat,n1393gat);
nor NOR2_241(n1476gat,n1858gat,n1590gat);
nor NOR3_191(n1407gat,n1393gat,n1409gat,n1677gat);
nor NOR3_192(n1412gat,n1411gat,n1406gat,n2981gat);
nor NOR3_193(n2663gat,n2586gat,n2660gat,n2307gat);
nor NOR2_242(n2662gat,n2660gat,n2586gat);
nor NOR2_243(n2238gat,n2448gat,n2444gat);
nor NOR3_194(n87gat,n743gat,n17gat,n293gat);
nor NOR2_244(n200gat,n199gat,n92gat);
nor NOR3_195(n184gat,n189gat,n188gat,n179gat);
nor NOR2_245(n196gat,n297gat,n195gat);
nor NOR2_246(n204gat,n200gat,n196gat);
nor NOR4_8(n2163gat,n1790gat,n1310gat,n2664gat,n2168gat);
nor NOR2_247(n2258gat,n2260gat,n2189gat);
nor NOR2_248(n2255gat,n2261gat,n2188gat);
nor NOR3_196(n2015gat,n2039gat,n1774gat,n1315gat);
nor NOR2_249(n2017gat,n1790gat,n2016gat);
nor NOR2_250(n2018gat,n2016gat,n2097gat);
nor NOR4_9(n2014gat,n2035gat,n2093gat,n2018gat,n2664gat);
nor NOR2_251(n2194gat,n2187gat,n1855gat);
nor NOR2_252(n2192gat,n2184gat,n1855gat);
nor NOR2_253(n2185gat,n2261gat,n2189gat);
nor NOR2_254(n2132gat,n2133gat,n2131gat);
nor NOR2_255(n2130gat,n2134gat,n2185gat);
nor NOR2_256(n2057gat,n2049gat,n1855gat);
nor NOR2_257(n2250gat,n2248gat,n2264gat);
nor NOR2_258(n2249gat,n2265gat,n3006gat);
nor NOR2_259(n2329gat,n1855gat,n3007gat);
nor NOR2_260(n1958gat,n1963gat,n1886gat);
nor NOR3_197(n1895gat,n1845gat,n1891gat,n1968gat);
nor NOR2_261(n1710gat,n1709gat,n1629gat);
nor NOR2_262(n1630gat,n1895gat,n1631gat);
nor NOR2_263(n2195gat,n2200gat,n1855gat);
nor NOR2_264(n2556gat,n1711gat,n2437gat);
nor NOR2_265(n2539gat,n2048gat,n2437gat);
nor NOR3_198(n1894gat,n1968gat,n1891gat,n1969gat);
nor NOR2_266(n1847gat,n1958gat,n1845gat);
nor NOR2_267(n1846gat,n1845gat,n1893gat);
nor NOR2_268(n2436gat,n2437gat,n1892gat);
nor NOR2_269(n2055gat,n1891gat,n1958gat);
nor NOR2_270(n1967gat,n1893gat,n1968gat);
nor NOR2_271(n2387gat,n2056gat,n2437gat);
nor NOR2_272(n1959gat,n1956gat,n1963gat);
nor NOR2_273(n1957gat,n1886gat,n1887gat);
nor NOR2_274(n2330gat,n2437gat,n1961gat);
nor NOR2_275(n2147gat,n2988gat,n1855gat);
nor NOR2_276(n2498gat,n2199gat,n2328gat);
nor NOR2_277(n2193gat,n2393gat,n2439gat);
nor NOR2_278(n2211gat,n2193gat,n2402gat);
nor NOR2_279(n2210gat,n2401gat,n2151gat);
nor NOR2_280(n2396gat,n2199gat,n2209gat);
nor NOR2_281(n2053gat,n2393gat,n2438gat);
nor NOR2_282(n1964gat,n2392gat,n2439gat);
nor NOR2_283(n2198gat,n2199gat,n2058gat);
nor NOR3_199(n2215gat,n2346gat,n2151gat,n2402gat);
nor NOR2_284(n2350gat,n2405gat,n2349gat);
nor NOR2_285(n2282gat,n2406gat,n2215gat);
nor NOR2_286(n2197gat,n2199gat,n2281gat);
nor NOR3_200(n2213gat,n2402gat,n2151gat,n2345gat);
nor NOR2_287(n2150gat,n2401gat,n2346gat);
nor NOR2_288(n2149gat,n2193gat,n2346gat);
nor NOR2_289(n2196gat,n2199gat,n2146gat);
nor NOR3_201(n1882gat,n2124gat,n2115gat,n2239gat);
nor NOR2_290(n1962gat,n1963gat,n1893gat);
nor NOR2_291(n1896gat,n2995gat,n1895gat);
nor NOR2_292(n1972gat,n1974gat,n1970gat);
nor NOR2_293(n1971gat,n1896gat,n1973gat);
nor NOR2_294(n2559gat,n2999gat,n2437gat);
nor NOR2_295(n2331gat,n2393gat,n2401gat);
nor NOR2_296(n2352gat,n3011gat,n2215gat);
nor NOR2_297(n2566gat,n2643gat,n2564gat);
nor NOR2_298(n2565gat,n2352gat,n2642gat);
nor NOR2_299(n2637gat,n3015gat,n2199gat);
nor NOR3_202(n84gat,n296gat,n17gat,n294gat);
nor NOR2_300(n89gat,n88gat,n2784gat);
nor NOR2_301(n110gat,n182gat,n89gat);
nor NOR2_302(n1074gat,n2775gat,n110gat);
nor NOR3_203(n141gat,n155gat,n253gat,n150gat);
nor NOR2_303(n38gat,n151gat,n233gat);
nor NOR2_304(n37gat,n151gat,n154gat);
nor NOR2_305(n872gat,n375gat,n800gat);
nor NOR2_306(n234gat,n155gat,n233gat);
nor NOR2_307(n137gat,n154gat,n253gat);
nor NOR2_308(n378gat,n375gat,n235gat);
nor NOR2_309(n377gat,n110gat,n2778gat);
nor NOR2_310(n869gat,n219gat,n2792gat);
nor NOR2_311(n212gat,n182gat,n78gat);
nor NOR3_204(n250gat,n329gat,n387gat,n334gat);
nor NOR2_312(n249gat,n386gat,n330gat);
nor NOR2_313(n248gat,n330gat,n1490gat);
nor NOR2_314(n453gat,n372gat,n452gat);
nor NOR2_315(n448gat,n111gat,n2846gat);
nor NOR2_316(n974gat,n2844gat,n111gat);
nor NOR2_317(n251gat,n1490gat,n387gat);
nor NOR2_318(n244gat,n334gat,n386gat);
nor NOR2_319(n973gat,n372gat,n333gat);
nor NOR2_320(n870gat,n2669gat,n219gat);
nor NOR2_321(n975gat,n111gat,n2852gat);
nor NOR3_205(n246gat,n330gat,n325gat,n334gat);
nor NOR2_322(n245gat,n386gat,n334gat);
nor NOR2_323(n460gat,n462gat,n2884gat);
nor NOR2_324(n459gat,n457gat,n461gat);
nor NOR2_325(n972gat,n372gat,n458gat);
nor NOR2_326(n969gat,n219gat,n2672gat);
nor NOR2_327(n971gat,n111gat,n2840gat);
nor NOR3_206(n247gat,n334gat,n387gat,n330gat);
nor NOR2_328(n145gat,n144gat,n325gat);
nor NOR2_329(n143gat,n326gat,n247gat);
nor NOR2_330(n970gat,n372gat,n878gat);
nor NOR2_331(n968gat,n2789gat,n219gat);
nor NOR2_332(n772gat,n111gat,n2842gat);
nor NOR3_207(n142gat,n382gat,n326gat,n144gat);
nor NOR2_333(n40gat,n325gat,n383gat);
nor NOR2_334(n39gat,n383gat,n247gat);
nor NOR2_335(n451gat,n134gat,n372gat);
nor NOR2_336(n446gat,n219gat,n2781gat);
nor NOR3_208(n139gat,n253gat,n151gat,n254gat);
nor NOR2_337(n136gat,n253gat,n154gat);
nor NOR2_338(n391gat,n252gat,n468gat);
nor NOR2_339(n390gat,n469gat,n2877gat);
nor NOR2_340(n1083gat,n381gat,n375gat);
nor NOR2_341(n1077gat,n110gat,n2672gat);
nor NOR3_209(n140gat,n151gat,n253gat,n155gat);
nor NOR2_342(n242gat,n254gat,n241gat);
nor NOR2_343(n240gat,n255gat,n140gat);
nor NOR2_344(n871gat,n802gat,n375gat);
nor NOR2_345(n797gat,n110gat,n2734gat);
nor NOR3_210(n324gat,n255gat,n146gat,n241gat);
nor NOR2_346(n238gat,n147gat,n254gat);
nor NOR2_347(n237gat,n140gat,n147gat);
nor NOR2_348(n1082gat,n375gat,n380gat);
nor NOR2_349(n796gat,n2731gat,n110gat);
nor NOR3_211(n85gat,n17gat,n294gat,n637gat);
nor NOR3_212(n180gat,n286gat,n188gat,n287gat);
nor NOR2_350(n68gat,n85gat,n180gat);
nor NOR3_213(n186gat,n189gat,n287gat,n288gat);
nor NOR2_351(n357gat,n2726gat,n2860gat);
nor NOR3_214(n82gat,n16gat,n295gat,n637gat);
nor NOR2_352(n12gat,n186gat,n82gat);
nor NOR2_353(n1599gat,n1691gat,n336gat);
nor NOR2_354(n1613gat,n1544gat,n1698gat);
nor NOR3_215(n1756gat,n2512gat,n1769gat,n1773gat);
nor NOR2_355(n1586gat,n1869gat,n1683gat);
nor NOR3_216(n1755gat,n1769gat,n1773gat,n2512gat);
nor NOR3_217(n2538gat,n2620gat,n2625gat,n2488gat);
nor NOR3_218(n2483gat,n2537gat,n2482gat,n2486gat);
nor NOR2_356(n1391gat,n1513gat,n2442gat);
nor NOR3_219(n1471gat,n1334gat,n1858gat,n1604gat);
nor NOR2_357(n1469gat,n1858gat,n1608gat);
nor NOR3_220(n1472gat,n1476gat,n1471gat,n1469gat);
nor NOR2_358(n1927gat,n1790gat,n1635gat);
nor NOR2_359(n1470gat,n1472gat,n1747gat);
nor NOR3_221(n1402gat,n1858gat,n1393gat,n1604gat);
nor NOR2_360(n1400gat,n1674gat,n1403gat);
nor NOR2_361(n1567gat,n1634gat,n1735gat);
nor NOR3_222(n1399gat,n1806gat,n1338gat,n1584gat);
nor NOR4_10(n1564gat,n1584gat,n1719gat,n1790gat,n1576gat);
nor NOR2_362(n1600gat,n1685gat,n1427gat);
nor NOR3_223(n1519gat,n1584gat,n1339gat,n1600gat);
nor NOR2_363(n1397gat,n1519gat,n1401gat);
nor NOR2_364(n1398gat,n1455gat,n1397gat);
nor NOR2_365(n2008gat,n2012gat,n1774gat);
nor NOR2_366(n2005gat,n2002gat,n2857gat);
nor NOR2_367(n1818gat,n1823gat,n2005gat);
nor NOR3_224(n1759gat,n1818gat,n1935gat,n2765gat);
nor NOR3_225(n1686gat,n1774gat,n1869gat,n1684gat);
nor NOR2_368(n1533gat,n1524gat,n1403gat);
nor NOR3_226(n1863gat,n1991gat,n2283gat,n1989gat);
nor NOR3_227(n1860gat,n1988gat,n2216gat,n1862gat);
nor NOR2_369(n1915gat,n1859gat,n1919gat);
nor NOR2_370(n1510gat,n1584gat,n1460gat);
nor NOR2_371(n1800gat,n1635gat,n1919gat);
nor NOR2_372(n1459gat,n1595gat,n1454gat);
nor NOR2_373(n1458gat,n1510gat,n1459gat);
nor NOR2_374(n1532gat,n1677gat,n1458gat);
nor NOR2_375(n1467gat,n2289gat,n1468gat);
nor NOR3_228(n1466gat,n1392gat,n1461gat,n1396gat);
nor NOR2_376(n1531gat,n1507gat,n1477gat);
nor NOR2_377(n1593gat,n1551gat,n1310gat);
nor NOR3_229(n1602gat,n1594gat,n1587gat,n2989gat);
nor NOR3_230(n1761gat,n2985gat,n1602gat,n1681gat);
nor NOR3_231(n1760gat,n1681gat,n1602gat,n2985gat);
nor NOR3_232(n1721gat,n2442gat,n1690gat,n1978gat);
nor NOR2_378(n520gat,n374gat,n2862gat);
nor NOR2_379(n519gat,n2854gat,n374gat);
nor NOR2_380(n518gat,n520gat,n519gat);
nor NOR2_381(n418gat,n374gat,n2723gat);
nor NOR2_382(n411gat,n374gat,n2726gat);
nor NOR2_383(n522gat,n374gat,n2859gat);
nor NOR2_384(n516gat,n374gat,n2715gat);
nor NOR4_11(n410gat,n417gat,n413gat,n412gat,n406gat);
nor NOR2_385(n354gat,n411gat,n522gat);
nor NOR3_233(n355gat,n517gat,n410gat,n354gat);
nor NOR2_386(n408gat,n516gat,n407gat);
nor NOR2_387(n526gat,n2859gat,n740gat);
nor NOR2_388(n531gat,n740gat,n2854gat);
nor NOR2_389(n530gat,n2862gat,n740gat);
nor NOR3_234(n525gat,n526gat,n531gat,n530gat);
nor NOR2_390(n356gat,n2726gat,n740gat);
nor NOR2_391(n415gat,n2723gat,n740gat);
nor NOR2_392(n521gat,n740gat,n2715gat);
nor NOR3_235(n532gat,n527gat,n416gat,n528gat);
nor NOR2_393(n359gat,n290gat,n358gat);
nor NOR2_394(n420gat,n408gat,n359gat);
nor NOR2_395(n523gat,n522gat,n356gat);
nor NOR2_396(n634gat,n418gat,n521gat);
nor NOR2_397(n414gat,n411gat,n415gat);
nor NOR3_236(n635gat,n639gat,n634gat,n414gat);
nor NOR2_398(n1100gat,n1297gat,n1111gat);
nor NOR3_237(n630gat,n634gat,n523gat,n524gat);
nor NOR2_399(n994gat,n1112gat,n882gat);
nor NOR3_238(n629gat,n414gat,n634gat,n523gat);
nor NOR2_400(n989gat,n721gat,n741gat);
nor NOR3_239(n632gat,n414gat,n523gat,n633gat);
nor NOR2_401(n880gat,n926gat,n566gat);
nor NOR3_240(n636gat,n414gat,n633gat,n639gat);
nor NOR2_402(n801gat,n672gat,n670gat);
nor NOR2_403(n879gat,n2931gat,n801gat);
nor NOR2_404(n1003gat,n420gat,n879gat);
nor NOR2_405(n1255gat,n1123gat,n1225gat);
nor NOR2_406(n1012gat,n1007gat,n918gat);
nor NOR2_407(n905gat,n625gat,n1006gat);
nor NOR2_408(n1009gat,n1255gat,n2943gat);
nor NOR2_409(n409gat,n406gat,n407gat);
nor NOR2_410(n292gat,n415gat,n356gat);
nor NOR2_411(n291gat,n290gat,n292gat);
nor NOR2_412(n419gat,n409gat,n291gat);
nor NOR2_413(n902gat,n1009gat,n419gat);
nor NOR2_414(n1099gat,n1111gat,n1293gat);
nor NOR2_415(n998gat,n725gat,n741gat);
nor NOR2_416(n995gat,n823gat,n1112gat);
nor NOR2_417(n980gat,n875gat,n926gat);
nor NOR2_418(n1001gat,n420gat,n1002gat);
nor NOR2_419(n1175gat,n621gat,n1006gat);
nor NOR2_420(n1174gat,n845gat,n1007gat);
nor NOR2_421(n1243gat,n1281gat,n1123gat);
nor NOR2_422(n1171gat,n2960gat,n1243gat);
nor NOR2_423(n999gat,n419gat,n1171gat);
nor NOR2_424(n1244gat,n1123gat,n1134gat);
nor NOR2_425(n1323gat,n1007gat,n401gat);
nor NOR2_426(n1264gat,n1006gat,n617gat);
nor NOR2_427(n1265gat,n1244gat,n2969gat);
nor NOR2_428(n892gat,n419gat,n1265gat);
nor NOR2_429(n981gat,n926gat,n873gat);
nor NOR2_430(n890gat,n741gat,n702gat);
nor NOR2_431(n889gat,n1111gat,n1079gat);
nor NOR2_432(n886gat,n683gat,n1112gat);
nor NOR2_433(n891gat,n420gat,n888gat);
nor NOR2_434(n904gat,n1006gat,n490gat);
nor NOR2_435(n903gat,n1007gat,n397gat);
nor NOR2_436(n1254gat,n1123gat,n1044gat);
nor NOR2_437(n1008gat,n2942gat,n1254gat);
nor NOR2_438(n900gat,n419gat,n1008gat);
nor NOR2_439(n1152gat,n926gat,n1150gat);
nor NOR2_440(n1092gat,n1147gat,n1111gat);
nor NOR2_441(n997gat,n741gat,n393gat);
nor NOR2_442(n993gat,n1112gat,n698gat);
nor NOR2_443(n895gat,n420gat,n898gat);
nor NOR2_444(n1094gat,n1112gat,n583gat);
nor NOR2_445(n1093gat,n1111gat,n864gat);
nor NOR2_446(n988gat,n340gat,n741gat);
nor NOR2_447(n984gat,n926gat,n983gat);
nor NOR2_448(n1178gat,n420gat,n1179gat);
nor NOR2_449(n1267gat,n613gat,n1006gat);
nor NOR2_450(n1257gat,n1007gat,n274gat);
nor NOR2_451(n1253gat,n930gat,n1123gat);
nor NOR2_452(n1266gat,n2965gat,n1253gat);
nor NOR2_453(n1116gat,n419gat,n1266gat);
nor NOR2_454(n1375gat,n1006gat,n706gat);
nor NOR2_455(n1324gat,n164gat,n1007gat);
nor NOR2_456(n1200gat,n1120gat,n1123gat);
nor NOR2_457(n1172gat,n2961gat,n1200gat);
nor NOR2_458(n899gat,n419gat,n1172gat);
nor NOR2_459(n1091gat,n1111gat,n956gat);
nor NOR2_460(n1088gat,n1085gat,n926gat);
nor NOR2_461(n992gat,n815gat,n1112gat);
nor NOR2_462(n987gat,n741gat,n159gat);
nor NOR2_463(n896gat,n897gat,n420gat);
nor NOR2_464(n1262gat,n837gat,n1006gat);
nor NOR2_465(n1260gat,n1007gat,n278gat);
nor NOR2_466(n1251gat,n1123gat,n1071gat);
nor NOR2_467(n1259gat,n2967gat,n1251gat);
nor NOR2_468(n901gat,n419gat,n1259gat);
nor NOR2_469(n1098gat,n336gat,n741gat);
nor NOR2_470(n1090gat,n1111gat,n860gat);
nor NOR2_471(n986gat,n985gat,n926gat);
nor NOR2_472(n885gat,n579gat,n1112gat);
nor NOR2_473(n893gat,n894gat,n420gat);
nor NOR2_474(n1097gat,n270gat,n741gat);
nor NOR2_475(n1089gat,n1067gat,n1111gat);
nor NOR2_476(n1087gat,n926gat,n1084gat);
nor NOR2_477(n991gat,n1112gat,n679gat);
nor NOR2_478(n1177gat,n1180gat,n420gat);
nor NOR2_479(n1212gat,n1123gat,n1034gat);
nor NOR2_480(n1326gat,n1007gat,n282gat);
nor NOR2_481(n1261gat,n833gat,n1006gat);
nor NOR2_482(n1263gat,n1212gat,n2968gat);
nor NOR2_483(n1115gat,n1263gat,n419gat);
nor NOR2_484(n977gat,n670gat,n671gat);
nor NOR3_241(n631gat,n523gat,n633gat,n524gat);
nor NOR2_485(n1096gat,n819gat,n1112gat);
nor NOR2_486(n1095gat,n1240gat,n1111gat);
nor NOR2_487(n990gat,n841gat,n741gat);
nor NOR2_488(n979gat,n1601gat,n926gat);
nor NOR2_489(n978gat,n2944gat,n2945gat);
nor NOR2_490(n1004gat,n978gat,n420gat);
nor NOR2_491(n1199gat,n1123gat,n1284gat);
nor NOR2_492(n1176gat,n829gat,n1006gat);
nor NOR2_493(n1173gat,n1007gat,n1025gat);
nor NOR2_494(n1252gat,n1199gat,n2962gat);
nor NOR2_495(n1000gat,n419gat,n1252gat);
nor NOR2_496(n1029gat,n978gat,n455gat);
nor NOR2_497(n1028gat,n455gat,n879gat);
nor NOR2_498(n1031gat,n1002gat,n455gat);
nor NOR2_499(n1030gat,n455gat,n888gat);
nor NOR2_500(n1011gat,n455gat,n898gat);
nor NOR2_501(n1181gat,n455gat,n1179gat);
nor NOR2_502(n1010gat,n897gat,n455gat);
nor NOR2_503(n1005gat,n894gat,n455gat);
nor NOR2_504(n1182gat,n1180gat,n455gat);
nor NOR2_505(n1757gat,n1773gat,n1769gat);
nor NOR2_506(n1745gat,n1869gat,n1757gat);
nor NOR2_507(n73gat,n67gat,n2784gat);
nor NOR2_508(n70gat,n71gat,n2720gat);
nor NOR2_509(n77gat,n76gat,n2784gat);
nor NOR2_510(n13gat,n2720gat,n14gat);

endmodule